module blk0(e0, out);
  input [4:0] e0;
  output [4:0] out;
  wire f;
  assign out[4:0] = 5'b01001;
endmodule
