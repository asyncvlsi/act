module blk0(e0, out);
  input [12:0] e0;
  output [12:0] out;
  wire f;
  assign out[12:0] = 13'b0100101110100;
endmodule
