module blk0(e0, out);
  input [4:0] e0;
  output [4:0] out;
  assign out = e0[4:0];
endmodule
