module blk_i0_4(out);
  (* src = "./exprop_0.v:12.7-12.13" *)
  wire _xtpa0;
  (* src = "./exprop_0.v:9.15-9.18" *)
  output [3:0] out;
  wire [3:0] out;
  assign _xtpa0 = 1'b0;
  assign out = 4'b0000;
endmodule
