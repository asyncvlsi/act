
module b14_DW01_add_7 ( A, B, CI, SUM, CO );
  input [30:1] A;
  input [30:0] B;
  output [30:0] SUM;
  input CI;
  output CO;
  wire   \A[2] , \A[1] , \A[0] , \carry[28] , \carry[27] , \carry[26] ,
         \carry[25] , \carry[24] , \carry[23] , \carry[22] , \carry[21] ,
         \carry[20] , \carry[19] , \carry[18] , \carry[17] , \carry[16] ,
         \carry[15] , \carry[14] , \carry[13] , \carry[12] , \carry[11] ,
         \carry[10] , \carry[9] , \carry[8] , \carry[7] , \carry[6] ,
         \carry[5] , \carry[4] ;
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign \carry[4]  = A[3];

  and2a3 U1 ( .A(A[28]), .B(\carry[28] ), .Y(SUM[29]) );
  xor2a1 U2 ( .A(A[28]), .B(\carry[28] ), .Y(SUM[28]) );
  and2a3 U3 ( .A(A[27]), .B(\carry[27] ), .Y(\carry[28] ) );
  xor2a1 U4 ( .A(A[27]), .B(\carry[27] ), .Y(SUM[27]) );
  and2a3 U5 ( .A(A[26]), .B(\carry[26] ), .Y(\carry[27] ) );
  xor2a1 U6 ( .A(A[26]), .B(\carry[26] ), .Y(SUM[26]) );
  and2a3 U7 ( .A(A[25]), .B(\carry[25] ), .Y(\carry[26] ) );
  xor2a1 U8 ( .A(A[25]), .B(\carry[25] ), .Y(SUM[25]) );
  and2a3 U9 ( .A(A[24]), .B(\carry[24] ), .Y(\carry[25] ) );
  xor2a1 U10 ( .A(A[24]), .B(\carry[24] ), .Y(SUM[24]) );
  and2a3 U11 ( .A(A[23]), .B(\carry[23] ), .Y(\carry[24] ) );
  xor2a1 U12 ( .A(A[23]), .B(\carry[23] ), .Y(SUM[23]) );
  and2a3 U13 ( .A(A[22]), .B(\carry[22] ), .Y(\carry[23] ) );
  xor2a1 U14 ( .A(A[22]), .B(\carry[22] ), .Y(SUM[22]) );
  and2a3 U15 ( .A(A[21]), .B(\carry[21] ), .Y(\carry[22] ) );
  xor2a1 U16 ( .A(A[21]), .B(\carry[21] ), .Y(SUM[21]) );
  and2a3 U17 ( .A(A[20]), .B(\carry[20] ), .Y(\carry[21] ) );
  xor2a1 U18 ( .A(A[20]), .B(\carry[20] ), .Y(SUM[20]) );
  and2a3 U19 ( .A(A[19]), .B(\carry[19] ), .Y(\carry[20] ) );
  xor2a1 U20 ( .A(A[19]), .B(\carry[19] ), .Y(SUM[19]) );
  and2a3 U21 ( .A(A[18]), .B(\carry[18] ), .Y(\carry[19] ) );
  xor2a1 U22 ( .A(A[18]), .B(\carry[18] ), .Y(SUM[18]) );
  and2a3 U23 ( .A(A[17]), .B(\carry[17] ), .Y(\carry[18] ) );
  xor2a1 U24 ( .A(A[17]), .B(\carry[17] ), .Y(SUM[17]) );
  and2a3 U25 ( .A(A[16]), .B(\carry[16] ), .Y(\carry[17] ) );
  xor2a1 U26 ( .A(A[16]), .B(\carry[16] ), .Y(SUM[16]) );
  and2a3 U27 ( .A(A[15]), .B(\carry[15] ), .Y(\carry[16] ) );
  xor2a1 U28 ( .A(A[15]), .B(\carry[15] ), .Y(SUM[15]) );
  and2a3 U29 ( .A(A[14]), .B(\carry[14] ), .Y(\carry[15] ) );
  xor2a1 U30 ( .A(A[14]), .B(\carry[14] ), .Y(SUM[14]) );
  and2a3 U31 ( .A(A[13]), .B(\carry[13] ), .Y(\carry[14] ) );
  xor2a1 U32 ( .A(A[13]), .B(\carry[13] ), .Y(SUM[13]) );
  and2a3 U33 ( .A(A[12]), .B(\carry[12] ), .Y(\carry[13] ) );
  xor2a1 U34 ( .A(A[12]), .B(\carry[12] ), .Y(SUM[12]) );
  and2a3 U35 ( .A(A[11]), .B(\carry[11] ), .Y(\carry[12] ) );
  xor2a1 U36 ( .A(A[11]), .B(\carry[11] ), .Y(SUM[11]) );
  and2a3 U37 ( .A(A[10]), .B(\carry[10] ), .Y(\carry[11] ) );
  xor2a1 U38 ( .A(A[10]), .B(\carry[10] ), .Y(SUM[10]) );
  and2a3 U39 ( .A(A[9]), .B(\carry[9] ), .Y(\carry[10] ) );
  xor2a1 U40 ( .A(A[9]), .B(\carry[9] ), .Y(SUM[9]) );
  and2a3 U41 ( .A(A[8]), .B(\carry[8] ), .Y(\carry[9] ) );
  xor2a1 U42 ( .A(A[8]), .B(\carry[8] ), .Y(SUM[8]) );
  and2a3 U43 ( .A(A[7]), .B(\carry[7] ), .Y(\carry[8] ) );
  xor2a1 U44 ( .A(A[7]), .B(\carry[7] ), .Y(SUM[7]) );
  and2a3 U45 ( .A(A[6]), .B(\carry[6] ), .Y(\carry[7] ) );
  xor2a1 U46 ( .A(A[6]), .B(\carry[6] ), .Y(SUM[6]) );
  and2a3 U47 ( .A(A[5]), .B(\carry[5] ), .Y(\carry[6] ) );
  xor2a1 U48 ( .A(A[5]), .B(\carry[5] ), .Y(SUM[5]) );
  and2a3 U49 ( .A(A[4]), .B(\carry[4] ), .Y(\carry[5] ) );
  xor2a1 U50 ( .A(A[4]), .B(\carry[4] ), .Y(SUM[4]) );
  inv1a1 U51 ( .A(\carry[4] ), .Y(SUM[3]) );
endmodule


module b14_DW01_sub_5 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , \carry[31] , \carry[30] , \carry[29] , \carry[28] ,
         \carry[27] , \carry[26] , \carry[25] , \carry[24] , \carry[23] ,
         \carry[22] , \carry[21] , \carry[20] , \carry[19] , \carry[18] ,
         \carry[17] , \carry[16] , \carry[15] , \carry[14] , \carry[13] ,
         \carry[12] , \carry[11] , \carry[10] , \carry[9] , \carry[8] ,
         \carry[7] , \carry[6] , \carry[5] , \carry[4] , \carry[3] ,
         \carry[2] , \carry[1] , \B_not[31] , \B_not[30] , \B_not[29] ,
         \B_not[28] , \B_not[27] , \B_not[26] , \B_not[25] , \B_not[24] ,
         \B_not[23] , \B_not[22] , \B_not[21] , \B_not[20] , \B_not[19] ,
         \B_not[18] , \B_not[17] , \B_not[16] , \B_not[15] , \B_not[14] ,
         \B_not[13] , \B_not[12] , \B_not[11] , \B_not[10] , \B_not[9] ,
         \B_not[8] , \B_not[7] , \B_not[6] , \B_not[5] , \B_not[4] ,
         \B_not[3] , \B_not[2] , \B_not[1] ;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  xor2a1 U1 ( .A(\B_not[31] ), .B(\carry[31] ), .Y(DIFF[31]) );
  and2a3 U2 ( .A(\B_not[30] ), .B(\carry[30] ), .Y(\carry[31] ) );
  xor2a1 U3 ( .A(\B_not[30] ), .B(\carry[30] ), .Y(DIFF[30]) );
  and2a3 U4 ( .A(\B_not[29] ), .B(\carry[29] ), .Y(\carry[30] ) );
  xor2a1 U5 ( .A(\B_not[29] ), .B(\carry[29] ), .Y(DIFF[29]) );
  and2a3 U6 ( .A(\B_not[28] ), .B(\carry[28] ), .Y(\carry[29] ) );
  xor2a1 U7 ( .A(\B_not[28] ), .B(\carry[28] ), .Y(DIFF[28]) );
  and2a3 U8 ( .A(\B_not[27] ), .B(\carry[27] ), .Y(\carry[28] ) );
  xor2a1 U9 ( .A(\B_not[27] ), .B(\carry[27] ), .Y(DIFF[27]) );
  and2a3 U10 ( .A(\B_not[26] ), .B(\carry[26] ), .Y(\carry[27] ) );
  xor2a1 U11 ( .A(\B_not[26] ), .B(\carry[26] ), .Y(DIFF[26]) );
  and2a3 U12 ( .A(\B_not[25] ), .B(\carry[25] ), .Y(\carry[26] ) );
  xor2a1 U13 ( .A(\B_not[25] ), .B(\carry[25] ), .Y(DIFF[25]) );
  and2a3 U14 ( .A(\B_not[24] ), .B(\carry[24] ), .Y(\carry[25] ) );
  xor2a1 U15 ( .A(\B_not[24] ), .B(\carry[24] ), .Y(DIFF[24]) );
  and2a3 U16 ( .A(\B_not[23] ), .B(\carry[23] ), .Y(\carry[24] ) );
  xor2a1 U17 ( .A(\B_not[23] ), .B(\carry[23] ), .Y(DIFF[23]) );
  and2a3 U18 ( .A(\B_not[22] ), .B(\carry[22] ), .Y(\carry[23] ) );
  xor2a1 U19 ( .A(\B_not[22] ), .B(\carry[22] ), .Y(DIFF[22]) );
  and2a3 U20 ( .A(\B_not[21] ), .B(\carry[21] ), .Y(\carry[22] ) );
  xor2a1 U21 ( .A(\B_not[21] ), .B(\carry[21] ), .Y(DIFF[21]) );
  and2a3 U22 ( .A(\B_not[20] ), .B(\carry[20] ), .Y(\carry[21] ) );
  xor2a1 U23 ( .A(\B_not[20] ), .B(\carry[20] ), .Y(DIFF[20]) );
  and2a3 U24 ( .A(\B_not[19] ), .B(\carry[19] ), .Y(\carry[20] ) );
  xor2a1 U25 ( .A(\B_not[19] ), .B(\carry[19] ), .Y(DIFF[19]) );
  and2a3 U26 ( .A(\B_not[18] ), .B(\carry[18] ), .Y(\carry[19] ) );
  xor2a1 U27 ( .A(\B_not[18] ), .B(\carry[18] ), .Y(DIFF[18]) );
  and2a3 U28 ( .A(\B_not[17] ), .B(\carry[17] ), .Y(\carry[18] ) );
  xor2a1 U29 ( .A(\B_not[17] ), .B(\carry[17] ), .Y(DIFF[17]) );
  and2a3 U30 ( .A(\B_not[16] ), .B(\carry[16] ), .Y(\carry[17] ) );
  xor2a1 U31 ( .A(\B_not[16] ), .B(\carry[16] ), .Y(DIFF[16]) );
  and2a3 U32 ( .A(\B_not[15] ), .B(\carry[15] ), .Y(\carry[16] ) );
  xor2a1 U33 ( .A(\B_not[15] ), .B(\carry[15] ), .Y(DIFF[15]) );
  and2a3 U34 ( .A(\B_not[14] ), .B(\carry[14] ), .Y(\carry[15] ) );
  xor2a1 U35 ( .A(\B_not[14] ), .B(\carry[14] ), .Y(DIFF[14]) );
  and2a3 U36 ( .A(\B_not[13] ), .B(\carry[13] ), .Y(\carry[14] ) );
  xor2a1 U37 ( .A(\B_not[13] ), .B(\carry[13] ), .Y(DIFF[13]) );
  and2a3 U38 ( .A(\B_not[12] ), .B(\carry[12] ), .Y(\carry[13] ) );
  xor2a1 U39 ( .A(\B_not[12] ), .B(\carry[12] ), .Y(DIFF[12]) );
  and2a3 U40 ( .A(\B_not[11] ), .B(\carry[11] ), .Y(\carry[12] ) );
  xor2a1 U41 ( .A(\B_not[11] ), .B(\carry[11] ), .Y(DIFF[11]) );
  and2a3 U42 ( .A(\B_not[10] ), .B(\carry[10] ), .Y(\carry[11] ) );
  xor2a1 U43 ( .A(\B_not[10] ), .B(\carry[10] ), .Y(DIFF[10]) );
  and2a3 U44 ( .A(\B_not[9] ), .B(\carry[9] ), .Y(\carry[10] ) );
  xor2a1 U45 ( .A(\B_not[9] ), .B(\carry[9] ), .Y(DIFF[9]) );
  and2a3 U46 ( .A(\B_not[8] ), .B(\carry[8] ), .Y(\carry[9] ) );
  xor2a1 U47 ( .A(\B_not[8] ), .B(\carry[8] ), .Y(DIFF[8]) );
  and2a3 U48 ( .A(\B_not[7] ), .B(\carry[7] ), .Y(\carry[8] ) );
  xor2a1 U49 ( .A(\B_not[7] ), .B(\carry[7] ), .Y(DIFF[7]) );
  and2a3 U50 ( .A(\B_not[6] ), .B(\carry[6] ), .Y(\carry[7] ) );
  xor2a1 U51 ( .A(\B_not[6] ), .B(\carry[6] ), .Y(DIFF[6]) );
  and2a3 U52 ( .A(\B_not[5] ), .B(\carry[5] ), .Y(\carry[6] ) );
  xor2a1 U53 ( .A(\B_not[5] ), .B(\carry[5] ), .Y(DIFF[5]) );
  and2a3 U54 ( .A(\B_not[4] ), .B(\carry[4] ), .Y(\carry[5] ) );
  xor2a1 U55 ( .A(\B_not[4] ), .B(\carry[4] ), .Y(DIFF[4]) );
  and2a3 U56 ( .A(\B_not[3] ), .B(\carry[3] ), .Y(\carry[4] ) );
  xor2a1 U57 ( .A(\B_not[3] ), .B(\carry[3] ), .Y(DIFF[3]) );
  and2a3 U58 ( .A(\B_not[2] ), .B(\carry[2] ), .Y(\carry[3] ) );
  xor2a1 U59 ( .A(\B_not[2] ), .B(\carry[2] ), .Y(DIFF[2]) );
  and2a3 U60 ( .A(\B_not[1] ), .B(\carry[1] ), .Y(\carry[2] ) );
  xor2a1 U61 ( .A(\B_not[1] ), .B(\carry[1] ), .Y(DIFF[1]) );
  inv1a1 U62 ( .A(\B[0] ), .Y(\carry[1] ) );
  inv1a1 U63 ( .A(B[9]), .Y(\B_not[9] ) );
  inv1a1 U64 ( .A(B[8]), .Y(\B_not[8] ) );
  inv1a1 U65 ( .A(B[7]), .Y(\B_not[7] ) );
  inv1a1 U66 ( .A(B[6]), .Y(\B_not[6] ) );
  inv1a1 U67 ( .A(B[5]), .Y(\B_not[5] ) );
  inv1a1 U68 ( .A(B[4]), .Y(\B_not[4] ) );
  inv1a1 U69 ( .A(B[3]), .Y(\B_not[3] ) );
  inv1a1 U70 ( .A(B[31]), .Y(\B_not[31] ) );
  inv1a1 U71 ( .A(B[30]), .Y(\B_not[30] ) );
  inv1a1 U72 ( .A(B[2]), .Y(\B_not[2] ) );
  inv1a1 U73 ( .A(B[29]), .Y(\B_not[29] ) );
  inv1a1 U74 ( .A(B[28]), .Y(\B_not[28] ) );
  inv1a1 U75 ( .A(B[27]), .Y(\B_not[27] ) );
  inv1a1 U76 ( .A(B[26]), .Y(\B_not[26] ) );
  inv1a1 U77 ( .A(B[25]), .Y(\B_not[25] ) );
  inv1a1 U78 ( .A(B[24]), .Y(\B_not[24] ) );
  inv1a1 U79 ( .A(B[23]), .Y(\B_not[23] ) );
  inv1a1 U80 ( .A(B[22]), .Y(\B_not[22] ) );
  inv1a1 U81 ( .A(B[21]), .Y(\B_not[21] ) );
  inv1a1 U82 ( .A(B[20]), .Y(\B_not[20] ) );
  inv1a1 U83 ( .A(B[1]), .Y(\B_not[1] ) );
  inv1a1 U84 ( .A(B[19]), .Y(\B_not[19] ) );
  inv1a1 U85 ( .A(B[18]), .Y(\B_not[18] ) );
  inv1a1 U86 ( .A(B[17]), .Y(\B_not[17] ) );
  inv1a1 U87 ( .A(B[16]), .Y(\B_not[16] ) );
  inv1a1 U88 ( .A(B[15]), .Y(\B_not[15] ) );
  inv1a1 U89 ( .A(B[14]), .Y(\B_not[14] ) );
  inv1a1 U90 ( .A(B[13]), .Y(\B_not[13] ) );
  inv1a1 U91 ( .A(B[12]), .Y(\B_not[12] ) );
  inv1a1 U92 ( .A(B[11]), .Y(\B_not[11] ) );
  inv1a1 U93 ( .A(B[10]), .Y(\B_not[10] ) );
endmodule


module b14_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , \carry[31] , \carry[30] , \carry[29] , \carry[28] ,
         \carry[27] , \carry[26] , \carry[25] , \carry[24] , \carry[23] ,
         \carry[22] , \carry[21] , \carry[20] , \carry[19] , \carry[18] ,
         \carry[17] , \carry[16] , \carry[15] , \carry[14] , \carry[13] ,
         \carry[12] , \carry[11] , \carry[10] , \carry[9] , \carry[8] ,
         \carry[7] , \carry[6] , \carry[5] , \carry[4] , \carry[3] ,
         \carry[2] , \carry[1] , \B_not[31] , \B_not[30] , \B_not[29] ,
         \B_not[28] , \B_not[27] , \B_not[26] , \B_not[25] , \B_not[24] ,
         \B_not[23] , \B_not[22] , \B_not[21] , \B_not[20] , \B_not[19] ,
         \B_not[18] , \B_not[17] , \B_not[16] , \B_not[15] , \B_not[14] ,
         \B_not[13] , \B_not[12] , \B_not[11] , \B_not[10] , \B_not[9] ,
         \B_not[8] , \B_not[7] , \B_not[6] , \B_not[5] , \B_not[4] ,
         \B_not[3] , \B_not[2] , \B_not[1] ;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  xor2a1 U1 ( .A(\B_not[31] ), .B(\carry[31] ), .Y(DIFF[31]) );
  and2a3 U2 ( .A(\B_not[30] ), .B(\carry[30] ), .Y(\carry[31] ) );
  xor2a1 U3 ( .A(\B_not[30] ), .B(\carry[30] ), .Y(DIFF[30]) );
  and2a3 U4 ( .A(\B_not[29] ), .B(\carry[29] ), .Y(\carry[30] ) );
  xor2a1 U5 ( .A(\B_not[29] ), .B(\carry[29] ), .Y(DIFF[29]) );
  and2a3 U6 ( .A(\B_not[28] ), .B(\carry[28] ), .Y(\carry[29] ) );
  xor2a1 U7 ( .A(\B_not[28] ), .B(\carry[28] ), .Y(DIFF[28]) );
  and2a3 U8 ( .A(\B_not[27] ), .B(\carry[27] ), .Y(\carry[28] ) );
  xor2a1 U9 ( .A(\B_not[27] ), .B(\carry[27] ), .Y(DIFF[27]) );
  and2a3 U10 ( .A(\B_not[26] ), .B(\carry[26] ), .Y(\carry[27] ) );
  xor2a1 U11 ( .A(\B_not[26] ), .B(\carry[26] ), .Y(DIFF[26]) );
  and2a3 U12 ( .A(\B_not[25] ), .B(\carry[25] ), .Y(\carry[26] ) );
  xor2a1 U13 ( .A(\B_not[25] ), .B(\carry[25] ), .Y(DIFF[25]) );
  and2a3 U14 ( .A(\B_not[24] ), .B(\carry[24] ), .Y(\carry[25] ) );
  xor2a1 U15 ( .A(\B_not[24] ), .B(\carry[24] ), .Y(DIFF[24]) );
  and2a3 U16 ( .A(\B_not[23] ), .B(\carry[23] ), .Y(\carry[24] ) );
  xor2a1 U17 ( .A(\B_not[23] ), .B(\carry[23] ), .Y(DIFF[23]) );
  and2a3 U18 ( .A(\B_not[22] ), .B(\carry[22] ), .Y(\carry[23] ) );
  xor2a1 U19 ( .A(\B_not[22] ), .B(\carry[22] ), .Y(DIFF[22]) );
  and2a3 U20 ( .A(\B_not[21] ), .B(\carry[21] ), .Y(\carry[22] ) );
  xor2a1 U21 ( .A(\B_not[21] ), .B(\carry[21] ), .Y(DIFF[21]) );
  and2a3 U22 ( .A(\B_not[20] ), .B(\carry[20] ), .Y(\carry[21] ) );
  xor2a1 U23 ( .A(\B_not[20] ), .B(\carry[20] ), .Y(DIFF[20]) );
  and2a3 U24 ( .A(\B_not[19] ), .B(\carry[19] ), .Y(\carry[20] ) );
  xor2a1 U25 ( .A(\B_not[19] ), .B(\carry[19] ), .Y(DIFF[19]) );
  and2a3 U26 ( .A(\B_not[18] ), .B(\carry[18] ), .Y(\carry[19] ) );
  xor2a1 U27 ( .A(\B_not[18] ), .B(\carry[18] ), .Y(DIFF[18]) );
  and2a3 U28 ( .A(\B_not[17] ), .B(\carry[17] ), .Y(\carry[18] ) );
  xor2a1 U29 ( .A(\B_not[17] ), .B(\carry[17] ), .Y(DIFF[17]) );
  and2a3 U30 ( .A(\B_not[16] ), .B(\carry[16] ), .Y(\carry[17] ) );
  xor2a1 U31 ( .A(\B_not[16] ), .B(\carry[16] ), .Y(DIFF[16]) );
  and2a3 U32 ( .A(\B_not[15] ), .B(\carry[15] ), .Y(\carry[16] ) );
  xor2a1 U33 ( .A(\B_not[15] ), .B(\carry[15] ), .Y(DIFF[15]) );
  and2a3 U34 ( .A(\B_not[14] ), .B(\carry[14] ), .Y(\carry[15] ) );
  xor2a1 U35 ( .A(\B_not[14] ), .B(\carry[14] ), .Y(DIFF[14]) );
  and2a3 U36 ( .A(\B_not[13] ), .B(\carry[13] ), .Y(\carry[14] ) );
  xor2a1 U37 ( .A(\B_not[13] ), .B(\carry[13] ), .Y(DIFF[13]) );
  and2a3 U38 ( .A(\B_not[12] ), .B(\carry[12] ), .Y(\carry[13] ) );
  xor2a1 U39 ( .A(\B_not[12] ), .B(\carry[12] ), .Y(DIFF[12]) );
  and2a3 U40 ( .A(\B_not[11] ), .B(\carry[11] ), .Y(\carry[12] ) );
  xor2a1 U41 ( .A(\B_not[11] ), .B(\carry[11] ), .Y(DIFF[11]) );
  and2a3 U42 ( .A(\B_not[10] ), .B(\carry[10] ), .Y(\carry[11] ) );
  xor2a1 U43 ( .A(\B_not[10] ), .B(\carry[10] ), .Y(DIFF[10]) );
  and2a3 U44 ( .A(\B_not[9] ), .B(\carry[9] ), .Y(\carry[10] ) );
  xor2a1 U45 ( .A(\B_not[9] ), .B(\carry[9] ), .Y(DIFF[9]) );
  and2a3 U46 ( .A(\B_not[8] ), .B(\carry[8] ), .Y(\carry[9] ) );
  xor2a1 U47 ( .A(\B_not[8] ), .B(\carry[8] ), .Y(DIFF[8]) );
  and2a3 U48 ( .A(\B_not[7] ), .B(\carry[7] ), .Y(\carry[8] ) );
  xor2a1 U49 ( .A(\B_not[7] ), .B(\carry[7] ), .Y(DIFF[7]) );
  and2a3 U50 ( .A(\B_not[6] ), .B(\carry[6] ), .Y(\carry[7] ) );
  xor2a1 U51 ( .A(\B_not[6] ), .B(\carry[6] ), .Y(DIFF[6]) );
  and2a3 U52 ( .A(\B_not[5] ), .B(\carry[5] ), .Y(\carry[6] ) );
  xor2a1 U53 ( .A(\B_not[5] ), .B(\carry[5] ), .Y(DIFF[5]) );
  and2a3 U54 ( .A(\B_not[4] ), .B(\carry[4] ), .Y(\carry[5] ) );
  xor2a1 U55 ( .A(\B_not[4] ), .B(\carry[4] ), .Y(DIFF[4]) );
  and2a3 U56 ( .A(\B_not[3] ), .B(\carry[3] ), .Y(\carry[4] ) );
  xor2a1 U57 ( .A(\B_not[3] ), .B(\carry[3] ), .Y(DIFF[3]) );
  and2a3 U58 ( .A(\B_not[2] ), .B(\carry[2] ), .Y(\carry[3] ) );
  xor2a1 U59 ( .A(\B_not[2] ), .B(\carry[2] ), .Y(DIFF[2]) );
  and2a3 U60 ( .A(\B_not[1] ), .B(\carry[1] ), .Y(\carry[2] ) );
  xor2a1 U61 ( .A(\B_not[1] ), .B(\carry[1] ), .Y(DIFF[1]) );
  inv1a1 U62 ( .A(\B[0] ), .Y(\carry[1] ) );
  inv1a1 U63 ( .A(B[9]), .Y(\B_not[9] ) );
  inv1a1 U64 ( .A(B[8]), .Y(\B_not[8] ) );
  inv1a1 U65 ( .A(B[7]), .Y(\B_not[7] ) );
  inv1a1 U66 ( .A(B[6]), .Y(\B_not[6] ) );
  inv1a1 U67 ( .A(B[5]), .Y(\B_not[5] ) );
  inv1a1 U68 ( .A(B[4]), .Y(\B_not[4] ) );
  inv1a1 U69 ( .A(B[3]), .Y(\B_not[3] ) );
  inv1a1 U70 ( .A(B[31]), .Y(\B_not[31] ) );
  inv1a1 U71 ( .A(B[30]), .Y(\B_not[30] ) );
  inv1a1 U72 ( .A(B[2]), .Y(\B_not[2] ) );
  inv1a1 U73 ( .A(B[29]), .Y(\B_not[29] ) );
  inv1a1 U74 ( .A(B[28]), .Y(\B_not[28] ) );
  inv1a1 U75 ( .A(B[27]), .Y(\B_not[27] ) );
  inv1a1 U76 ( .A(B[26]), .Y(\B_not[26] ) );
  inv1a1 U77 ( .A(B[25]), .Y(\B_not[25] ) );
  inv1a1 U78 ( .A(B[24]), .Y(\B_not[24] ) );
  inv1a1 U79 ( .A(B[23]), .Y(\B_not[23] ) );
  inv1a1 U80 ( .A(B[22]), .Y(\B_not[22] ) );
  inv1a1 U81 ( .A(B[21]), .Y(\B_not[21] ) );
  inv1a1 U82 ( .A(B[20]), .Y(\B_not[20] ) );
  inv1a1 U83 ( .A(B[1]), .Y(\B_not[1] ) );
  inv1a1 U84 ( .A(B[19]), .Y(\B_not[19] ) );
  inv1a1 U85 ( .A(B[18]), .Y(\B_not[18] ) );
  inv1a1 U86 ( .A(B[17]), .Y(\B_not[17] ) );
  inv1a1 U87 ( .A(B[16]), .Y(\B_not[16] ) );
  inv1a1 U88 ( .A(B[15]), .Y(\B_not[15] ) );
  inv1a1 U89 ( .A(B[14]), .Y(\B_not[14] ) );
  inv1a1 U90 ( .A(B[13]), .Y(\B_not[13] ) );
  inv1a1 U91 ( .A(B[12]), .Y(\B_not[12] ) );
  inv1a1 U92 ( .A(B[11]), .Y(\B_not[11] ) );
  inv1a1 U93 ( .A(B[10]), .Y(\B_not[10] ) );
endmodule


module b14_DW01_add_5 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   \carry[19] , \carry[18] , \carry[17] , \carry[16] , \carry[15] ,
         \carry[14] , \carry[13] , \carry[12] , \carry[11] , \carry[10] ,
         \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] , \carry[2] , \carry[1] ;

  xor3a1 U1_19 ( .A(A[19]), .B(B[19]), .C(\carry[19] ), .Y(SUM[19]) );
  fa1a1 U1_13 ( .A(A[13]), .B(B[13]), .CI(\carry[13] ), .CO(\carry[14] ), .S(
        SUM[13]) );
  fa1a1 U1_11 ( .A(A[11]), .B(B[11]), .CI(\carry[11] ), .CO(\carry[12] ), .S(
        SUM[11]) );
  fa1a1 U1_9 ( .A(A[9]), .B(B[9]), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  fa1a1 U1_7 ( .A(A[7]), .B(B[7]), .CI(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  fa1a1 U1_5 ( .A(A[5]), .B(B[5]), .CI(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  fa1a1 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  fa1a1 U1_1 ( .A(A[1]), .B(B[1]), .CI(\carry[1] ), .CO(\carry[2] ), .S(SUM[1]) );
  fa1a1 U1_6 ( .A(A[6]), .B(B[6]), .CI(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  fa1a1 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  fa1a1 U1_10 ( .A(A[10]), .B(B[10]), .CI(\carry[10] ), .CO(\carry[11] ), .S(
        SUM[10]) );
  fa1a1 U1_12 ( .A(A[12]), .B(B[12]), .CI(\carry[12] ), .CO(\carry[13] ), .S(
        SUM[12]) );
  fa1a1 U1_14 ( .A(A[14]), .B(B[14]), .CI(\carry[14] ), .CO(\carry[15] ), .S(
        SUM[14]) );
  fa1a1 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  fa1a1 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  fa1a1 U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), .S(
        SUM[17]) );
  fa1a1 U1_15 ( .A(A[15]), .B(B[15]), .CI(\carry[15] ), .CO(\carry[16] ), .S(
        SUM[15]) );
  fa1a1 U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  fa1a1 U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  and2a3 U1 ( .A(B[0]), .B(A[0]), .Y(\carry[1] ) );
  xor2a1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module b14_DW01_add_4 ( A, B, CI, SUM, CO );
  input [19:0] A;
  input [19:0] B;
  output [19:0] SUM;
  input CI;
  output CO;
  wire   \carry[19] , \carry[18] , \carry[17] , \carry[16] , \carry[15] ,
         \carry[14] , \carry[13] , \carry[12] , \carry[11] , \carry[10] ,
         \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] , \carry[2] , \carry[1] ;

  xor3a1 U1_19 ( .A(A[19]), .B(B[19]), .C(\carry[19] ), .Y(SUM[19]) );
  fa1a1 U1_13 ( .A(A[13]), .B(B[13]), .CI(\carry[13] ), .CO(\carry[14] ), .S(
        SUM[13]) );
  fa1a1 U1_11 ( .A(A[11]), .B(B[11]), .CI(\carry[11] ), .CO(\carry[12] ), .S(
        SUM[11]) );
  fa1a1 U1_9 ( .A(A[9]), .B(B[9]), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  fa1a1 U1_7 ( .A(A[7]), .B(B[7]), .CI(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  fa1a1 U1_5 ( .A(A[5]), .B(B[5]), .CI(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  fa1a1 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  fa1a1 U1_1 ( .A(A[1]), .B(B[1]), .CI(\carry[1] ), .CO(\carry[2] ), .S(SUM[1]) );
  fa1a1 U1_6 ( .A(A[6]), .B(B[6]), .CI(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  fa1a1 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  fa1a1 U1_10 ( .A(A[10]), .B(B[10]), .CI(\carry[10] ), .CO(\carry[11] ), .S(
        SUM[10]) );
  fa1a1 U1_12 ( .A(A[12]), .B(B[12]), .CI(\carry[12] ), .CO(\carry[13] ), .S(
        SUM[12]) );
  fa1a1 U1_14 ( .A(A[14]), .B(B[14]), .CI(\carry[14] ), .CO(\carry[15] ), .S(
        SUM[14]) );
  fa1a1 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  fa1a1 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  fa1a1 U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), .S(
        SUM[17]) );
  fa1a1 U1_15 ( .A(A[15]), .B(B[15]), .CI(\carry[15] ), .CO(\carry[16] ), .S(
        SUM[15]) );
  fa1a1 U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  fa1a1 U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  and2a3 U1 ( .A(B[0]), .B(A[0]), .Y(\carry[1] ) );
  xor2a1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module b14_DW01_add_3 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   \carry[29] , \carry[28] , \carry[27] , \carry[26] , \carry[25] ,
         \carry[24] , \carry[23] , \carry[22] , \carry[21] , \carry[20] ,
         \carry[19] , \carry[18] , \carry[17] , \carry[16] , \carry[15] ,
         \carry[14] , \carry[13] , \carry[12] , \carry[11] , \carry[10] ,
         \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] , \carry[2] , \carry[1] ;

  xor3a3 U1_29 ( .A(A[29]), .B(B[29]), .C(\carry[29] ), .Y(SUM[29]) );
  fa1a1 U1_27 ( .A(A[27]), .B(B[27]), .CI(\carry[27] ), .CO(\carry[28] ), .S(
        SUM[27]) );
  fa1a1 U1_23 ( .A(A[23]), .B(B[23]), .CI(\carry[23] ), .CO(\carry[24] ), .S(
        SUM[23]) );
  fa1a1 U1_22 ( .A(A[22]), .B(B[22]), .CI(\carry[22] ), .CO(\carry[23] ), .S(
        SUM[22]) );
  fa1a1 U1_26 ( .A(A[26]), .B(B[26]), .CI(\carry[26] ), .CO(\carry[27] ), .S(
        SUM[26]) );
  fa1a1 U1_28 ( .A(A[28]), .B(B[28]), .CI(\carry[28] ), .CO(\carry[29] ), .S(
        SUM[28]) );
  fa1a1 U1_25 ( .A(A[25]), .B(B[25]), .CI(\carry[25] ), .CO(\carry[26] ), .S(
        SUM[25]) );
  fa1a1 U1_21 ( .A(A[21]), .B(B[21]), .CI(\carry[21] ), .CO(\carry[22] ), .S(
        SUM[21]) );
  fa1a1 U1_20 ( .A(A[20]), .B(B[20]), .CI(\carry[20] ), .CO(\carry[21] ), .S(
        SUM[20]) );
  fa1a1 U1_24 ( .A(A[24]), .B(B[24]), .CI(\carry[24] ), .CO(\carry[25] ), .S(
        SUM[24]) );
  fa1a1 U1_19 ( .A(A[19]), .B(B[19]), .CI(\carry[19] ), .CO(\carry[20] ), .S(
        SUM[19]) );
  fa1a1 U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), .S(
        SUM[17]) );
  fa1a1 U1_13 ( .A(A[13]), .B(B[13]), .CI(\carry[13] ), .CO(\carry[14] ), .S(
        SUM[13]) );
  fa1a1 U1_9 ( .A(A[9]), .B(B[9]), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  fa1a1 U1_5 ( .A(A[5]), .B(B[5]), .CI(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  fa1a1 U1_1 ( .A(A[1]), .B(B[1]), .CI(\carry[1] ), .CO(\carry[2] ), .S(SUM[1]) );
  fa1a1 U1_15 ( .A(A[15]), .B(B[15]), .CI(\carry[15] ), .CO(\carry[16] ), .S(
        SUM[15]) );
  fa1a1 U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  fa1a1 U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  fa1a1 U1_11 ( .A(A[11]), .B(B[11]), .CI(\carry[11] ), .CO(\carry[12] ), .S(
        SUM[11]) );
  fa1a1 U1_7 ( .A(A[7]), .B(B[7]), .CI(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  fa1a1 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  fa1a1 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  fa1a1 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  fa1a1 U1_6 ( .A(A[6]), .B(B[6]), .CI(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  fa1a1 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  fa1a1 U1_10 ( .A(A[10]), .B(B[10]), .CI(\carry[10] ), .CO(\carry[11] ), .S(
        SUM[10]) );
  fa1a1 U1_12 ( .A(A[12]), .B(B[12]), .CI(\carry[12] ), .CO(\carry[13] ), .S(
        SUM[12]) );
  fa1a1 U1_14 ( .A(A[14]), .B(B[14]), .CI(\carry[14] ), .CO(\carry[15] ), .S(
        SUM[14]) );
  and2a3 U1 ( .A(B[0]), .B(A[0]), .Y(\carry[1] ) );
  xor2a1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module b14_DW01_add_2 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   \carry[29] , \carry[28] , \carry[27] , \carry[26] , \carry[25] ,
         \carry[24] , \carry[23] , \carry[22] , \carry[21] , \carry[20] ,
         \carry[19] , \carry[18] , \carry[17] , \carry[16] , \carry[15] ,
         \carry[14] , \carry[13] , \carry[12] , \carry[11] , \carry[10] ,
         \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] , \carry[2] , \carry[1] ;

  fa1a1 U1_28 ( .A(A[28]), .B(B[28]), .CI(\carry[28] ), .CO(\carry[29] ), .S(
        SUM[28]) );
  fa1a1 U1_27 ( .A(A[27]), .B(B[27]), .CI(\carry[27] ), .CO(\carry[28] ), .S(
        SUM[27]) );
  fa1a1 U1_26 ( .A(A[26]), .B(B[26]), .CI(\carry[26] ), .CO(\carry[27] ), .S(
        SUM[26]) );
  fa1a1 U1_23 ( .A(A[23]), .B(B[23]), .CI(\carry[23] ), .CO(\carry[24] ), .S(
        SUM[23]) );
  fa1a1 U1_22 ( .A(A[22]), .B(B[22]), .CI(\carry[22] ), .CO(\carry[23] ), .S(
        SUM[22]) );
  fa1a1 U1_25 ( .A(A[25]), .B(B[25]), .CI(\carry[25] ), .CO(\carry[26] ), .S(
        SUM[25]) );
  fa1a1 U1_24 ( .A(A[24]), .B(B[24]), .CI(\carry[24] ), .CO(\carry[25] ), .S(
        SUM[24]) );
  fa1a1 U1_21 ( .A(A[21]), .B(B[21]), .CI(\carry[21] ), .CO(\carry[22] ), .S(
        SUM[21]) );
  fa1a1 U1_20 ( .A(A[20]), .B(B[20]), .CI(\carry[20] ), .CO(\carry[21] ), .S(
        SUM[20]) );
  xor3a3 U1_29 ( .A(A[29]), .B(B[29]), .C(\carry[29] ), .Y(SUM[29]) );
  fa1a1 U1_19 ( .A(A[19]), .B(B[19]), .CI(\carry[19] ), .CO(\carry[20] ), .S(
        SUM[19]) );
  fa1a1 U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), .S(
        SUM[17]) );
  fa1a1 U1_13 ( .A(A[13]), .B(B[13]), .CI(\carry[13] ), .CO(\carry[14] ), .S(
        SUM[13]) );
  fa1a1 U1_9 ( .A(A[9]), .B(B[9]), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  fa1a1 U1_5 ( .A(A[5]), .B(B[5]), .CI(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  fa1a1 U1_1 ( .A(A[1]), .B(B[1]), .CI(\carry[1] ), .CO(\carry[2] ), .S(SUM[1]) );
  fa1a1 U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  fa1a1 U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  fa1a1 U1_15 ( .A(A[15]), .B(B[15]), .CI(\carry[15] ), .CO(\carry[16] ), .S(
        SUM[15]) );
  fa1a1 U1_14 ( .A(A[14]), .B(B[14]), .CI(\carry[14] ), .CO(\carry[15] ), .S(
        SUM[14]) );
  fa1a1 U1_12 ( .A(A[12]), .B(B[12]), .CI(\carry[12] ), .CO(\carry[13] ), .S(
        SUM[12]) );
  fa1a1 U1_11 ( .A(A[11]), .B(B[11]), .CI(\carry[11] ), .CO(\carry[12] ), .S(
        SUM[11]) );
  fa1a1 U1_10 ( .A(A[10]), .B(B[10]), .CI(\carry[10] ), .CO(\carry[11] ), .S(
        SUM[10]) );
  fa1a1 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  fa1a1 U1_7 ( .A(A[7]), .B(B[7]), .CI(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  fa1a1 U1_6 ( .A(A[6]), .B(B[6]), .CI(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  fa1a1 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  fa1a1 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  fa1a1 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  and2a3 U1 ( .A(B[0]), .B(A[0]), .Y(\carry[1] ) );
  xor2a1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module b14_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] DIFF;
  input CI;
  output CO;
  wire   \carry[29] , \carry[28] , \carry[27] , \carry[26] , \carry[25] ,
         \carry[24] , \carry[23] , \carry[22] , \carry[21] , \carry[20] ,
         \carry[19] , \carry[18] , \carry[17] , \carry[16] , \carry[15] ,
         \carry[14] , \carry[13] , \carry[12] , \carry[11] , \carry[10] ,
         \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] , \carry[2] , \carry[1] , \B_not[29] ,
         \B_not[28] , \B_not[27] , \B_not[26] , \B_not[25] , \B_not[24] ,
         \B_not[23] , \B_not[22] , \B_not[21] , \B_not[20] , \B_not[19] ,
         \B_not[18] , \B_not[17] , \B_not[16] , \B_not[15] , \B_not[14] ,
         \B_not[13] , \B_not[12] , \B_not[11] , \B_not[10] , \B_not[9] ,
         \B_not[8] , \B_not[7] , \B_not[6] , \B_not[5] , \B_not[4] ,
         \B_not[3] , \B_not[2] , \B_not[1] , \B_not[0] , n1;

  fa1a1 U2_28 ( .A(A[28]), .B(\B_not[28] ), .CI(\carry[28] ), .CO(\carry[29] ), 
        .S(DIFF[28]) );
  fa1a1 U2_27 ( .A(A[27]), .B(\B_not[27] ), .CI(\carry[27] ), .CO(\carry[28] ), 
        .S(DIFF[27]) );
  fa1a1 U2_26 ( .A(A[26]), .B(\B_not[26] ), .CI(\carry[26] ), .CO(\carry[27] ), 
        .S(DIFF[26]) );
  fa1a1 U2_23 ( .A(A[23]), .B(\B_not[23] ), .CI(\carry[23] ), .CO(\carry[24] ), 
        .S(DIFF[23]) );
  fa1a1 U2_22 ( .A(A[22]), .B(\B_not[22] ), .CI(\carry[22] ), .CO(\carry[23] ), 
        .S(DIFF[22]) );
  fa1a1 U2_19 ( .A(A[19]), .B(\B_not[19] ), .CI(\carry[19] ), .CO(\carry[20] ), 
        .S(DIFF[19]) );
  fa1a1 U2_25 ( .A(A[25]), .B(\B_not[25] ), .CI(\carry[25] ), .CO(\carry[26] ), 
        .S(DIFF[25]) );
  fa1a1 U2_24 ( .A(A[24]), .B(\B_not[24] ), .CI(\carry[24] ), .CO(\carry[25] ), 
        .S(DIFF[24]) );
  fa1a1 U2_21 ( .A(A[21]), .B(\B_not[21] ), .CI(\carry[21] ), .CO(\carry[22] ), 
        .S(DIFF[21]) );
  fa1a1 U2_20 ( .A(A[20]), .B(\B_not[20] ), .CI(\carry[20] ), .CO(\carry[21] ), 
        .S(DIFF[20]) );
  fa1a1 U2_18 ( .A(A[18]), .B(\B_not[18] ), .CI(\carry[18] ), .CO(\carry[19] ), 
        .S(DIFF[18]) );
  fa1a1 U2_15 ( .A(A[15]), .B(\B_not[15] ), .CI(\carry[15] ), .CO(\carry[16] ), 
        .S(DIFF[15]) );
  fa1a1 U2_14 ( .A(A[14]), .B(\B_not[14] ), .CI(\carry[14] ), .CO(\carry[15] ), 
        .S(DIFF[14]) );
  fa1a1 U2_11 ( .A(A[11]), .B(\B_not[11] ), .CI(\carry[11] ), .CO(\carry[12] ), 
        .S(DIFF[11]) );
  fa1a1 U2_10 ( .A(A[10]), .B(\B_not[10] ), .CI(\carry[10] ), .CO(\carry[11] ), 
        .S(DIFF[10]) );
  fa1a1 U2_7 ( .A(A[7]), .B(\B_not[7] ), .CI(\carry[7] ), .CO(\carry[8] ), .S(
        DIFF[7]) );
  fa1a1 U2_6 ( .A(A[6]), .B(\B_not[6] ), .CI(\carry[6] ), .CO(\carry[7] ), .S(
        DIFF[6]) );
  fa1a1 U2_3 ( .A(A[3]), .B(\B_not[3] ), .CI(\carry[3] ), .CO(\carry[4] ), .S(
        DIFF[3]) );
  fa1a1 U2_2 ( .A(A[2]), .B(\B_not[2] ), .CI(\carry[2] ), .CO(\carry[3] ), .S(
        DIFF[2]) );
  fa1a1 U2_17 ( .A(A[17]), .B(\B_not[17] ), .CI(\carry[17] ), .CO(\carry[18] ), 
        .S(DIFF[17]) );
  fa1a1 U2_16 ( .A(A[16]), .B(\B_not[16] ), .CI(\carry[16] ), .CO(\carry[17] ), 
        .S(DIFF[16]) );
  fa1a1 U2_13 ( .A(A[13]), .B(\B_not[13] ), .CI(\carry[13] ), .CO(\carry[14] ), 
        .S(DIFF[13]) );
  fa1a1 U2_12 ( .A(A[12]), .B(\B_not[12] ), .CI(\carry[12] ), .CO(\carry[13] ), 
        .S(DIFF[12]) );
  fa1a1 U2_9 ( .A(A[9]), .B(\B_not[9] ), .CI(\carry[9] ), .CO(\carry[10] ), 
        .S(DIFF[9]) );
  fa1a1 U2_8 ( .A(A[8]), .B(\B_not[8] ), .CI(\carry[8] ), .CO(\carry[9] ), .S(
        DIFF[8]) );
  fa1a1 U2_5 ( .A(A[5]), .B(\B_not[5] ), .CI(\carry[5] ), .CO(\carry[6] ), .S(
        DIFF[5]) );
  fa1a1 U2_4 ( .A(A[4]), .B(\B_not[4] ), .CI(\carry[4] ), .CO(\carry[5] ), .S(
        DIFF[4]) );
  fa1a1 U2_1 ( .A(A[1]), .B(\B_not[1] ), .CI(\carry[1] ), .CO(\carry[2] ), .S(
        DIFF[1]) );
  xor3a3 U2_29 ( .A(A[29]), .B(\B_not[29] ), .C(\carry[29] ), .Y(DIFF[29]) );
  or2a1 U1 ( .A(A[0]), .B(\B_not[0] ), .Y(\carry[1] ) );
  xor2a1 U2 ( .A(n1), .B(\B_not[0] ), .Y(DIFF[0]) );
  inv1a1 U3 ( .A(A[0]), .Y(n1) );
  inv1a1 U4 ( .A(B[9]), .Y(\B_not[9] ) );
  inv1a1 U5 ( .A(B[8]), .Y(\B_not[8] ) );
  inv1a1 U6 ( .A(B[7]), .Y(\B_not[7] ) );
  inv1a1 U7 ( .A(B[6]), .Y(\B_not[6] ) );
  inv1a1 U8 ( .A(B[5]), .Y(\B_not[5] ) );
  inv1a1 U9 ( .A(B[4]), .Y(\B_not[4] ) );
  inv1a1 U10 ( .A(B[3]), .Y(\B_not[3] ) );
  inv1a1 U11 ( .A(B[2]), .Y(\B_not[2] ) );
  inv1a1 U12 ( .A(B[29]), .Y(\B_not[29] ) );
  inv1a1 U13 ( .A(B[28]), .Y(\B_not[28] ) );
  inv1a1 U14 ( .A(B[27]), .Y(\B_not[27] ) );
  inv1a1 U15 ( .A(B[26]), .Y(\B_not[26] ) );
  inv1a1 U16 ( .A(B[25]), .Y(\B_not[25] ) );
  inv1a1 U17 ( .A(B[24]), .Y(\B_not[24] ) );
  inv1a1 U18 ( .A(B[23]), .Y(\B_not[23] ) );
  inv1a1 U19 ( .A(B[22]), .Y(\B_not[22] ) );
  inv1a1 U20 ( .A(B[21]), .Y(\B_not[21] ) );
  inv1a1 U21 ( .A(B[20]), .Y(\B_not[20] ) );
  inv1a1 U22 ( .A(B[1]), .Y(\B_not[1] ) );
  inv1a1 U23 ( .A(B[19]), .Y(\B_not[19] ) );
  inv1a1 U24 ( .A(B[18]), .Y(\B_not[18] ) );
  inv1a1 U25 ( .A(B[17]), .Y(\B_not[17] ) );
  inv1a1 U26 ( .A(B[16]), .Y(\B_not[16] ) );
  inv1a1 U27 ( .A(B[15]), .Y(\B_not[15] ) );
  inv1a1 U28 ( .A(B[14]), .Y(\B_not[14] ) );
  inv1a1 U29 ( .A(B[13]), .Y(\B_not[13] ) );
  inv1a1 U30 ( .A(B[12]), .Y(\B_not[12] ) );
  inv1a1 U31 ( .A(B[11]), .Y(\B_not[11] ) );
  inv1a1 U32 ( .A(B[10]), .Y(\B_not[10] ) );
  inv1a1 U33 ( .A(B[0]), .Y(\B_not[0] ) );
endmodule


module b14_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] DIFF;
  input CI;
  output CO;
  wire   \carry[29] , \carry[28] , \carry[27] , \carry[26] , \carry[25] ,
         \carry[24] , \carry[23] , \carry[22] , \carry[21] , \carry[20] ,
         \carry[19] , \carry[18] , \carry[17] , \carry[16] , \carry[15] ,
         \carry[14] , \carry[13] , \carry[12] , \carry[11] , \carry[10] ,
         \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] , \carry[2] , \carry[1] , \B_not[29] ,
         \B_not[28] , \B_not[27] , \B_not[26] , \B_not[25] , \B_not[24] ,
         \B_not[23] , \B_not[22] , \B_not[21] , \B_not[20] , \B_not[19] ,
         \B_not[18] , \B_not[17] , \B_not[16] , \B_not[15] , \B_not[14] ,
         \B_not[13] , \B_not[12] , \B_not[11] , \B_not[10] , \B_not[9] ,
         \B_not[8] , \B_not[7] , \B_not[6] , \B_not[5] , \B_not[4] ,
         \B_not[3] , \B_not[2] , \B_not[1] , \B_not[0] , n1;

  xor3a3 U2_29 ( .A(A[29]), .B(\B_not[29] ), .C(\carry[29] ), .Y(DIFF[29]) );
  fa1a1 U2_27 ( .A(A[27]), .B(\B_not[27] ), .CI(\carry[27] ), .CO(\carry[28] ), 
        .S(DIFF[27]) );
  fa1a1 U2_23 ( .A(A[23]), .B(\B_not[23] ), .CI(\carry[23] ), .CO(\carry[24] ), 
        .S(DIFF[23]) );
  fa1a1 U2_22 ( .A(A[22]), .B(\B_not[22] ), .CI(\carry[22] ), .CO(\carry[23] ), 
        .S(DIFF[22]) );
  fa1a1 U2_26 ( .A(A[26]), .B(\B_not[26] ), .CI(\carry[26] ), .CO(\carry[27] ), 
        .S(DIFF[26]) );
  fa1a1 U2_28 ( .A(A[28]), .B(\B_not[28] ), .CI(\carry[28] ), .CO(\carry[29] ), 
        .S(DIFF[28]) );
  fa1a1 U2_19 ( .A(A[19]), .B(\B_not[19] ), .CI(\carry[19] ), .CO(\carry[20] ), 
        .S(DIFF[19]) );
  fa1a1 U2_25 ( .A(A[25]), .B(\B_not[25] ), .CI(\carry[25] ), .CO(\carry[26] ), 
        .S(DIFF[25]) );
  fa1a1 U2_21 ( .A(A[21]), .B(\B_not[21] ), .CI(\carry[21] ), .CO(\carry[22] ), 
        .S(DIFF[21]) );
  fa1a1 U2_20 ( .A(A[20]), .B(\B_not[20] ), .CI(\carry[20] ), .CO(\carry[21] ), 
        .S(DIFF[20]) );
  fa1a1 U2_24 ( .A(A[24]), .B(\B_not[24] ), .CI(\carry[24] ), .CO(\carry[25] ), 
        .S(DIFF[24]) );
  fa1a1 U2_15 ( .A(A[15]), .B(\B_not[15] ), .CI(\carry[15] ), .CO(\carry[16] ), 
        .S(DIFF[15]) );
  fa1a1 U2_11 ( .A(A[11]), .B(\B_not[11] ), .CI(\carry[11] ), .CO(\carry[12] ), 
        .S(DIFF[11]) );
  fa1a1 U2_7 ( .A(A[7]), .B(\B_not[7] ), .CI(\carry[7] ), .CO(\carry[8] ), .S(
        DIFF[7]) );
  fa1a1 U2_3 ( .A(A[3]), .B(\B_not[3] ), .CI(\carry[3] ), .CO(\carry[4] ), .S(
        DIFF[3]) );
  fa1a1 U2_2 ( .A(A[2]), .B(\B_not[2] ), .CI(\carry[2] ), .CO(\carry[3] ), .S(
        DIFF[2]) );
  fa1a1 U2_6 ( .A(A[6]), .B(\B_not[6] ), .CI(\carry[6] ), .CO(\carry[7] ), .S(
        DIFF[6]) );
  fa1a1 U2_10 ( .A(A[10]), .B(\B_not[10] ), .CI(\carry[10] ), .CO(\carry[11] ), 
        .S(DIFF[10]) );
  fa1a1 U2_14 ( .A(A[14]), .B(\B_not[14] ), .CI(\carry[14] ), .CO(\carry[15] ), 
        .S(DIFF[14]) );
  fa1a1 U2_18 ( .A(A[18]), .B(\B_not[18] ), .CI(\carry[18] ), .CO(\carry[19] ), 
        .S(DIFF[18]) );
  fa1a1 U2_17 ( .A(A[17]), .B(\B_not[17] ), .CI(\carry[17] ), .CO(\carry[18] ), 
        .S(DIFF[17]) );
  fa1a1 U2_13 ( .A(A[13]), .B(\B_not[13] ), .CI(\carry[13] ), .CO(\carry[14] ), 
        .S(DIFF[13]) );
  fa1a1 U2_9 ( .A(A[9]), .B(\B_not[9] ), .CI(\carry[9] ), .CO(\carry[10] ), 
        .S(DIFF[9]) );
  fa1a1 U2_5 ( .A(A[5]), .B(\B_not[5] ), .CI(\carry[5] ), .CO(\carry[6] ), .S(
        DIFF[5]) );
  fa1a1 U2_4 ( .A(A[4]), .B(\B_not[4] ), .CI(\carry[4] ), .CO(\carry[5] ), .S(
        DIFF[4]) );
  fa1a1 U2_8 ( .A(A[8]), .B(\B_not[8] ), .CI(\carry[8] ), .CO(\carry[9] ), .S(
        DIFF[8]) );
  fa1a1 U2_12 ( .A(A[12]), .B(\B_not[12] ), .CI(\carry[12] ), .CO(\carry[13] ), 
        .S(DIFF[12]) );
  fa1a1 U2_16 ( .A(A[16]), .B(\B_not[16] ), .CI(\carry[16] ), .CO(\carry[17] ), 
        .S(DIFF[16]) );
  fa1a1 U2_1 ( .A(A[1]), .B(\B_not[1] ), .CI(\carry[1] ), .CO(\carry[2] ), .S(
        DIFF[1]) );
  or2a1 U1 ( .A(A[0]), .B(\B_not[0] ), .Y(\carry[1] ) );
  xor2a1 U2 ( .A(n1), .B(\B_not[0] ), .Y(DIFF[0]) );
  inv1a1 U3 ( .A(A[0]), .Y(n1) );
  inv1a1 U4 ( .A(B[9]), .Y(\B_not[9] ) );
  inv1a1 U5 ( .A(B[8]), .Y(\B_not[8] ) );
  inv1a1 U6 ( .A(B[7]), .Y(\B_not[7] ) );
  inv1a1 U7 ( .A(B[6]), .Y(\B_not[6] ) );
  inv1a1 U8 ( .A(B[5]), .Y(\B_not[5] ) );
  inv1a1 U9 ( .A(B[4]), .Y(\B_not[4] ) );
  inv1a1 U10 ( .A(B[3]), .Y(\B_not[3] ) );
  inv1a1 U11 ( .A(B[2]), .Y(\B_not[2] ) );
  inv1a1 U12 ( .A(B[29]), .Y(\B_not[29] ) );
  inv1a1 U13 ( .A(B[28]), .Y(\B_not[28] ) );
  inv1a1 U14 ( .A(B[27]), .Y(\B_not[27] ) );
  inv1a1 U15 ( .A(B[26]), .Y(\B_not[26] ) );
  inv1a1 U16 ( .A(B[25]), .Y(\B_not[25] ) );
  inv1a1 U17 ( .A(B[24]), .Y(\B_not[24] ) );
  inv1a1 U18 ( .A(B[23]), .Y(\B_not[23] ) );
  inv1a1 U19 ( .A(B[22]), .Y(\B_not[22] ) );
  inv1a1 U20 ( .A(B[21]), .Y(\B_not[21] ) );
  inv1a1 U21 ( .A(B[20]), .Y(\B_not[20] ) );
  inv1a1 U22 ( .A(B[1]), .Y(\B_not[1] ) );
  inv1a1 U23 ( .A(B[19]), .Y(\B_not[19] ) );
  inv1a1 U24 ( .A(B[18]), .Y(\B_not[18] ) );
  inv1a1 U25 ( .A(B[17]), .Y(\B_not[17] ) );
  inv1a1 U26 ( .A(B[16]), .Y(\B_not[16] ) );
  inv1a1 U27 ( .A(B[15]), .Y(\B_not[15] ) );
  inv1a1 U28 ( .A(B[14]), .Y(\B_not[14] ) );
  inv1a1 U29 ( .A(B[13]), .Y(\B_not[13] ) );
  inv1a1 U30 ( .A(B[12]), .Y(\B_not[12] ) );
  inv1a1 U31 ( .A(B[11]), .Y(\B_not[11] ) );
  inv1a1 U32 ( .A(B[10]), .Y(\B_not[10] ) );
  inv1a1 U33 ( .A(B[0]), .Y(\B_not[0] ) );
endmodule


module b14_DW01_add_1 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   \carry[29] , \carry[28] , \carry[27] , \carry[26] , \carry[25] ,
         \carry[24] , \carry[23] , \carry[22] , \carry[21] , \carry[20] ,
         \carry[19] , \carry[18] , \carry[17] , \carry[16] , \carry[15] ,
         \carry[14] , \carry[13] , \carry[12] , \carry[11] , \carry[10] ,
         \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] , \carry[2] , \carry[1] ;

  fa1a1 U1_28 ( .A(A[28]), .B(B[28]), .CI(\carry[28] ), .CO(\carry[29] ), .S(
        SUM[28]) );
  fa1a1 U1_27 ( .A(A[27]), .B(B[27]), .CI(\carry[27] ), .CO(\carry[28] ), .S(
        SUM[27]) );
  fa1a1 U1_26 ( .A(A[26]), .B(B[26]), .CI(\carry[26] ), .CO(\carry[27] ), .S(
        SUM[26]) );
  fa1a1 U1_23 ( .A(A[23]), .B(B[23]), .CI(\carry[23] ), .CO(\carry[24] ), .S(
        SUM[23]) );
  fa1a1 U1_22 ( .A(A[22]), .B(B[22]), .CI(\carry[22] ), .CO(\carry[23] ), .S(
        SUM[22]) );
  fa1a1 U1_25 ( .A(A[25]), .B(B[25]), .CI(\carry[25] ), .CO(\carry[26] ), .S(
        SUM[25]) );
  fa1a1 U1_24 ( .A(A[24]), .B(B[24]), .CI(\carry[24] ), .CO(\carry[25] ), .S(
        SUM[24]) );
  fa1a1 U1_21 ( .A(A[21]), .B(B[21]), .CI(\carry[21] ), .CO(\carry[22] ), .S(
        SUM[21]) );
  fa1a1 U1_20 ( .A(A[20]), .B(B[20]), .CI(\carry[20] ), .CO(\carry[21] ), .S(
        SUM[20]) );
  fa1a1 U1_19 ( .A(A[19]), .B(B[19]), .CI(\carry[19] ), .CO(\carry[20] ), .S(
        SUM[19]) );
  fa1a1 U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), .S(
        SUM[17]) );
  fa1a1 U1_13 ( .A(A[13]), .B(B[13]), .CI(\carry[13] ), .CO(\carry[14] ), .S(
        SUM[13]) );
  fa1a1 U1_9 ( .A(A[9]), .B(B[9]), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  fa1a1 U1_5 ( .A(A[5]), .B(B[5]), .CI(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  fa1a1 U1_1 ( .A(A[1]), .B(B[1]), .CI(\carry[1] ), .CO(\carry[2] ), .S(SUM[1]) );
  fa1a1 U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  fa1a1 U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  fa1a1 U1_15 ( .A(A[15]), .B(B[15]), .CI(\carry[15] ), .CO(\carry[16] ), .S(
        SUM[15]) );
  fa1a1 U1_14 ( .A(A[14]), .B(B[14]), .CI(\carry[14] ), .CO(\carry[15] ), .S(
        SUM[14]) );
  fa1a1 U1_12 ( .A(A[12]), .B(B[12]), .CI(\carry[12] ), .CO(\carry[13] ), .S(
        SUM[12]) );
  fa1a1 U1_11 ( .A(A[11]), .B(B[11]), .CI(\carry[11] ), .CO(\carry[12] ), .S(
        SUM[11]) );
  fa1a1 U1_10 ( .A(A[10]), .B(B[10]), .CI(\carry[10] ), .CO(\carry[11] ), .S(
        SUM[10]) );
  fa1a1 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  fa1a1 U1_7 ( .A(A[7]), .B(B[7]), .CI(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  fa1a1 U1_6 ( .A(A[6]), .B(B[6]), .CI(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  fa1a1 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  fa1a1 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  fa1a1 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  xor3a3 U1_29 ( .A(A[29]), .B(B[29]), .C(\carry[29] ), .Y(SUM[29]) );
  and2a3 U1 ( .A(B[0]), .B(A[0]), .Y(\carry[1] ) );
  xor2a1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module b14_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] DIFF;
  input CI;
  output CO;
  wire   \carry[29] , \carry[28] , \carry[27] , \carry[26] , \carry[25] ,
         \carry[24] , \carry[23] , \carry[22] , \carry[21] , \carry[20] ,
         \carry[19] , \carry[18] , \carry[17] , \carry[16] , \carry[15] ,
         \carry[14] , \carry[13] , \carry[12] , \carry[11] , \carry[10] ,
         \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] , \carry[2] , \carry[1] , \B_not[29] ,
         \B_not[28] , \B_not[27] , \B_not[26] , \B_not[25] , \B_not[24] ,
         \B_not[23] , \B_not[22] , \B_not[21] , \B_not[20] , \B_not[19] ,
         \B_not[18] , \B_not[17] , \B_not[16] , \B_not[15] , \B_not[14] ,
         \B_not[13] , \B_not[12] , \B_not[11] , \B_not[10] , \B_not[9] ,
         \B_not[8] , \B_not[7] , \B_not[6] , \B_not[5] , \B_not[4] ,
         \B_not[3] , \B_not[2] , \B_not[1] , \B_not[0] , n1;

  fa1a1 U2_28 ( .A(A[28]), .B(\B_not[28] ), .CI(\carry[28] ), .CO(\carry[29] ), 
        .S(DIFF[28]) );
  fa1a1 U2_27 ( .A(A[27]), .B(\B_not[27] ), .CI(\carry[27] ), .CO(\carry[28] ), 
        .S(DIFF[27]) );
  fa1a1 U2_26 ( .A(A[26]), .B(\B_not[26] ), .CI(\carry[26] ), .CO(\carry[27] ), 
        .S(DIFF[26]) );
  fa1a1 U2_23 ( .A(A[23]), .B(\B_not[23] ), .CI(\carry[23] ), .CO(\carry[24] ), 
        .S(DIFF[23]) );
  fa1a1 U2_22 ( .A(A[22]), .B(\B_not[22] ), .CI(\carry[22] ), .CO(\carry[23] ), 
        .S(DIFF[22]) );
  fa1a1 U2_19 ( .A(A[19]), .B(\B_not[19] ), .CI(\carry[19] ), .CO(\carry[20] ), 
        .S(DIFF[19]) );
  fa1a1 U2_25 ( .A(A[25]), .B(\B_not[25] ), .CI(\carry[25] ), .CO(\carry[26] ), 
        .S(DIFF[25]) );
  fa1a1 U2_24 ( .A(A[24]), .B(\B_not[24] ), .CI(\carry[24] ), .CO(\carry[25] ), 
        .S(DIFF[24]) );
  fa1a1 U2_21 ( .A(A[21]), .B(\B_not[21] ), .CI(\carry[21] ), .CO(\carry[22] ), 
        .S(DIFF[21]) );
  fa1a1 U2_20 ( .A(A[20]), .B(\B_not[20] ), .CI(\carry[20] ), .CO(\carry[21] ), 
        .S(DIFF[20]) );
  fa1a1 U2_18 ( .A(A[18]), .B(\B_not[18] ), .CI(\carry[18] ), .CO(\carry[19] ), 
        .S(DIFF[18]) );
  fa1a1 U2_15 ( .A(A[15]), .B(\B_not[15] ), .CI(\carry[15] ), .CO(\carry[16] ), 
        .S(DIFF[15]) );
  fa1a1 U2_14 ( .A(A[14]), .B(\B_not[14] ), .CI(\carry[14] ), .CO(\carry[15] ), 
        .S(DIFF[14]) );
  fa1a1 U2_11 ( .A(A[11]), .B(\B_not[11] ), .CI(\carry[11] ), .CO(\carry[12] ), 
        .S(DIFF[11]) );
  fa1a1 U2_10 ( .A(A[10]), .B(\B_not[10] ), .CI(\carry[10] ), .CO(\carry[11] ), 
        .S(DIFF[10]) );
  fa1a1 U2_7 ( .A(A[7]), .B(\B_not[7] ), .CI(\carry[7] ), .CO(\carry[8] ), .S(
        DIFF[7]) );
  fa1a1 U2_6 ( .A(A[6]), .B(\B_not[6] ), .CI(\carry[6] ), .CO(\carry[7] ), .S(
        DIFF[6]) );
  fa1a1 U2_3 ( .A(A[3]), .B(\B_not[3] ), .CI(\carry[3] ), .CO(\carry[4] ), .S(
        DIFF[3]) );
  fa1a1 U2_2 ( .A(A[2]), .B(\B_not[2] ), .CI(\carry[2] ), .CO(\carry[3] ), .S(
        DIFF[2]) );
  fa1a1 U2_17 ( .A(A[17]), .B(\B_not[17] ), .CI(\carry[17] ), .CO(\carry[18] ), 
        .S(DIFF[17]) );
  fa1a1 U2_16 ( .A(A[16]), .B(\B_not[16] ), .CI(\carry[16] ), .CO(\carry[17] ), 
        .S(DIFF[16]) );
  fa1a1 U2_13 ( .A(A[13]), .B(\B_not[13] ), .CI(\carry[13] ), .CO(\carry[14] ), 
        .S(DIFF[13]) );
  fa1a1 U2_12 ( .A(A[12]), .B(\B_not[12] ), .CI(\carry[12] ), .CO(\carry[13] ), 
        .S(DIFF[12]) );
  fa1a1 U2_9 ( .A(A[9]), .B(\B_not[9] ), .CI(\carry[9] ), .CO(\carry[10] ), 
        .S(DIFF[9]) );
  fa1a1 U2_8 ( .A(A[8]), .B(\B_not[8] ), .CI(\carry[8] ), .CO(\carry[9] ), .S(
        DIFF[8]) );
  fa1a1 U2_5 ( .A(A[5]), .B(\B_not[5] ), .CI(\carry[5] ), .CO(\carry[6] ), .S(
        DIFF[5]) );
  fa1a1 U2_4 ( .A(A[4]), .B(\B_not[4] ), .CI(\carry[4] ), .CO(\carry[5] ), .S(
        DIFF[4]) );
  fa1a1 U2_1 ( .A(A[1]), .B(\B_not[1] ), .CI(\carry[1] ), .CO(\carry[2] ), .S(
        DIFF[1]) );
  xor3a3 U2_29 ( .A(A[29]), .B(\B_not[29] ), .C(\carry[29] ), .Y(DIFF[29]) );
  or2a1 U1 ( .A(A[0]), .B(\B_not[0] ), .Y(\carry[1] ) );
  xor2a1 U2 ( .A(n1), .B(\B_not[0] ), .Y(DIFF[0]) );
  inv1a1 U3 ( .A(A[0]), .Y(n1) );
  inv1a1 U4 ( .A(B[9]), .Y(\B_not[9] ) );
  inv1a1 U5 ( .A(B[8]), .Y(\B_not[8] ) );
  inv1a1 U6 ( .A(B[7]), .Y(\B_not[7] ) );
  inv1a1 U7 ( .A(B[6]), .Y(\B_not[6] ) );
  inv1a1 U8 ( .A(B[5]), .Y(\B_not[5] ) );
  inv1a1 U9 ( .A(B[4]), .Y(\B_not[4] ) );
  inv1a1 U10 ( .A(B[3]), .Y(\B_not[3] ) );
  inv1a1 U11 ( .A(B[2]), .Y(\B_not[2] ) );
  inv1a1 U12 ( .A(B[29]), .Y(\B_not[29] ) );
  inv1a1 U13 ( .A(B[28]), .Y(\B_not[28] ) );
  inv1a1 U14 ( .A(B[27]), .Y(\B_not[27] ) );
  inv1a1 U15 ( .A(B[26]), .Y(\B_not[26] ) );
  inv1a1 U16 ( .A(B[25]), .Y(\B_not[25] ) );
  inv1a1 U17 ( .A(B[24]), .Y(\B_not[24] ) );
  inv1a1 U18 ( .A(B[23]), .Y(\B_not[23] ) );
  inv1a1 U19 ( .A(B[22]), .Y(\B_not[22] ) );
  inv1a1 U20 ( .A(B[21]), .Y(\B_not[21] ) );
  inv1a1 U21 ( .A(B[20]), .Y(\B_not[20] ) );
  inv1a1 U22 ( .A(B[1]), .Y(\B_not[1] ) );
  inv1a1 U23 ( .A(B[19]), .Y(\B_not[19] ) );
  inv1a1 U24 ( .A(B[18]), .Y(\B_not[18] ) );
  inv1a1 U25 ( .A(B[17]), .Y(\B_not[17] ) );
  inv1a1 U26 ( .A(B[16]), .Y(\B_not[16] ) );
  inv1a1 U27 ( .A(B[15]), .Y(\B_not[15] ) );
  inv1a1 U28 ( .A(B[14]), .Y(\B_not[14] ) );
  inv1a1 U29 ( .A(B[13]), .Y(\B_not[13] ) );
  inv1a1 U30 ( .A(B[12]), .Y(\B_not[12] ) );
  inv1a1 U31 ( .A(B[11]), .Y(\B_not[11] ) );
  inv1a1 U32 ( .A(B[10]), .Y(\B_not[10] ) );
  inv1a1 U33 ( .A(B[0]), .Y(\B_not[0] ) );
endmodule


module b14_DW01_add_0 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   \carry[29] , \carry[28] , \carry[27] , \carry[26] , \carry[25] ,
         \carry[24] , \carry[23] , \carry[22] , \carry[21] , \carry[20] ,
         \carry[19] , \carry[18] , \carry[17] , \carry[16] , \carry[15] ,
         \carry[14] , \carry[13] , \carry[12] , \carry[11] , \carry[10] ,
         \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] , \carry[2] , \carry[1] ;

  fa1a1 U1_28 ( .A(A[28]), .B(B[28]), .CI(\carry[28] ), .CO(\carry[29] ), .S(
        SUM[28]) );
  fa1a1 U1_27 ( .A(A[27]), .B(B[27]), .CI(\carry[27] ), .CO(\carry[28] ), .S(
        SUM[27]) );
  fa1a1 U1_26 ( .A(A[26]), .B(B[26]), .CI(\carry[26] ), .CO(\carry[27] ), .S(
        SUM[26]) );
  fa1a1 U1_23 ( .A(A[23]), .B(B[23]), .CI(\carry[23] ), .CO(\carry[24] ), .S(
        SUM[23]) );
  fa1a1 U1_22 ( .A(A[22]), .B(B[22]), .CI(\carry[22] ), .CO(\carry[23] ), .S(
        SUM[22]) );
  fa1a1 U1_25 ( .A(A[25]), .B(B[25]), .CI(\carry[25] ), .CO(\carry[26] ), .S(
        SUM[25]) );
  fa1a1 U1_24 ( .A(A[24]), .B(B[24]), .CI(\carry[24] ), .CO(\carry[25] ), .S(
        SUM[24]) );
  fa1a1 U1_21 ( .A(A[21]), .B(B[21]), .CI(\carry[21] ), .CO(\carry[22] ), .S(
        SUM[21]) );
  fa1a1 U1_20 ( .A(A[20]), .B(B[20]), .CI(\carry[20] ), .CO(\carry[21] ), .S(
        SUM[20]) );
  xor3a3 U1_29 ( .A(A[29]), .B(B[29]), .C(\carry[29] ), .Y(SUM[29]) );
  fa1a1 U1_19 ( .A(A[19]), .B(B[19]), .CI(\carry[19] ), .CO(\carry[20] ), .S(
        SUM[19]) );
  fa1a1 U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), .S(
        SUM[17]) );
  fa1a1 U1_13 ( .A(A[13]), .B(B[13]), .CI(\carry[13] ), .CO(\carry[14] ), .S(
        SUM[13]) );
  fa1a1 U1_9 ( .A(A[9]), .B(B[9]), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  fa1a1 U1_5 ( .A(A[5]), .B(B[5]), .CI(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  fa1a1 U1_1 ( .A(A[1]), .B(B[1]), .CI(\carry[1] ), .CO(\carry[2] ), .S(SUM[1]) );
  fa1a1 U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  fa1a1 U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  fa1a1 U1_15 ( .A(A[15]), .B(B[15]), .CI(\carry[15] ), .CO(\carry[16] ), .S(
        SUM[15]) );
  fa1a1 U1_14 ( .A(A[14]), .B(B[14]), .CI(\carry[14] ), .CO(\carry[15] ), .S(
        SUM[14]) );
  fa1a1 U1_12 ( .A(A[12]), .B(B[12]), .CI(\carry[12] ), .CO(\carry[13] ), .S(
        SUM[12]) );
  fa1a1 U1_11 ( .A(A[11]), .B(B[11]), .CI(\carry[11] ), .CO(\carry[12] ), .S(
        SUM[11]) );
  fa1a1 U1_10 ( .A(A[10]), .B(B[10]), .CI(\carry[10] ), .CO(\carry[11] ), .S(
        SUM[10]) );
  fa1a1 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  fa1a1 U1_7 ( .A(A[7]), .B(B[7]), .CI(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  fa1a1 U1_6 ( .A(A[6]), .B(B[6]), .CI(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  fa1a1 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  fa1a1 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  fa1a1 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  and2a3 U1 ( .A(B[0]), .B(A[0]), .Y(\carry[1] ) );
  xor2a1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module b14_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] DIFF;
  input CI;
  output CO;
  wire   \carry[29] , \carry[28] , \carry[27] , \carry[26] , \carry[25] ,
         \carry[24] , \carry[23] , \carry[22] , \carry[21] , \carry[20] ,
         \carry[19] , \carry[18] , \carry[17] , \carry[16] , \carry[15] ,
         \carry[14] , \carry[13] , \carry[12] , \carry[11] , \carry[10] ,
         \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] , \carry[2] , \carry[1] , \B_not[29] ,
         \B_not[28] , \B_not[27] , \B_not[26] , \B_not[25] , \B_not[24] ,
         \B_not[23] , \B_not[22] , \B_not[21] , \B_not[20] , \B_not[19] ,
         \B_not[18] , \B_not[17] , \B_not[16] , \B_not[15] , \B_not[14] ,
         \B_not[13] , \B_not[12] , \B_not[11] , \B_not[10] , \B_not[9] ,
         \B_not[8] , \B_not[7] , \B_not[6] , \B_not[5] , \B_not[4] ,
         \B_not[3] , \B_not[2] , \B_not[1] , \B_not[0] , n1;

  fa1a1 U2_28 ( .A(A[28]), .B(\B_not[28] ), .CI(\carry[28] ), .CO(\carry[29] ), 
        .S(DIFF[28]) );
  fa1a1 U2_27 ( .A(A[27]), .B(\B_not[27] ), .CI(\carry[27] ), .CO(\carry[28] ), 
        .S(DIFF[27]) );
  fa1a1 U2_26 ( .A(A[26]), .B(\B_not[26] ), .CI(\carry[26] ), .CO(\carry[27] ), 
        .S(DIFF[26]) );
  fa1a1 U2_23 ( .A(A[23]), .B(\B_not[23] ), .CI(\carry[23] ), .CO(\carry[24] ), 
        .S(DIFF[23]) );
  fa1a1 U2_22 ( .A(A[22]), .B(\B_not[22] ), .CI(\carry[22] ), .CO(\carry[23] ), 
        .S(DIFF[22]) );
  fa1a1 U2_19 ( .A(A[19]), .B(\B_not[19] ), .CI(\carry[19] ), .CO(\carry[20] ), 
        .S(DIFF[19]) );
  fa1a1 U2_25 ( .A(A[25]), .B(\B_not[25] ), .CI(\carry[25] ), .CO(\carry[26] ), 
        .S(DIFF[25]) );
  fa1a1 U2_24 ( .A(A[24]), .B(\B_not[24] ), .CI(\carry[24] ), .CO(\carry[25] ), 
        .S(DIFF[24]) );
  fa1a1 U2_21 ( .A(A[21]), .B(\B_not[21] ), .CI(\carry[21] ), .CO(\carry[22] ), 
        .S(DIFF[21]) );
  fa1a1 U2_20 ( .A(A[20]), .B(\B_not[20] ), .CI(\carry[20] ), .CO(\carry[21] ), 
        .S(DIFF[20]) );
  fa1a1 U2_18 ( .A(A[18]), .B(\B_not[18] ), .CI(\carry[18] ), .CO(\carry[19] ), 
        .S(DIFF[18]) );
  fa1a1 U2_15 ( .A(A[15]), .B(\B_not[15] ), .CI(\carry[15] ), .CO(\carry[16] ), 
        .S(DIFF[15]) );
  fa1a1 U2_14 ( .A(A[14]), .B(\B_not[14] ), .CI(\carry[14] ), .CO(\carry[15] ), 
        .S(DIFF[14]) );
  fa1a1 U2_11 ( .A(A[11]), .B(\B_not[11] ), .CI(\carry[11] ), .CO(\carry[12] ), 
        .S(DIFF[11]) );
  fa1a1 U2_10 ( .A(A[10]), .B(\B_not[10] ), .CI(\carry[10] ), .CO(\carry[11] ), 
        .S(DIFF[10]) );
  fa1a1 U2_7 ( .A(A[7]), .B(\B_not[7] ), .CI(\carry[7] ), .CO(\carry[8] ), .S(
        DIFF[7]) );
  fa1a1 U2_6 ( .A(A[6]), .B(\B_not[6] ), .CI(\carry[6] ), .CO(\carry[7] ), .S(
        DIFF[6]) );
  fa1a1 U2_3 ( .A(A[3]), .B(\B_not[3] ), .CI(\carry[3] ), .CO(\carry[4] ), .S(
        DIFF[3]) );
  fa1a1 U2_2 ( .A(A[2]), .B(\B_not[2] ), .CI(\carry[2] ), .CO(\carry[3] ), .S(
        DIFF[2]) );
  fa1a1 U2_17 ( .A(A[17]), .B(\B_not[17] ), .CI(\carry[17] ), .CO(\carry[18] ), 
        .S(DIFF[17]) );
  fa1a1 U2_16 ( .A(A[16]), .B(\B_not[16] ), .CI(\carry[16] ), .CO(\carry[17] ), 
        .S(DIFF[16]) );
  fa1a1 U2_13 ( .A(A[13]), .B(\B_not[13] ), .CI(\carry[13] ), .CO(\carry[14] ), 
        .S(DIFF[13]) );
  fa1a1 U2_12 ( .A(A[12]), .B(\B_not[12] ), .CI(\carry[12] ), .CO(\carry[13] ), 
        .S(DIFF[12]) );
  fa1a1 U2_9 ( .A(A[9]), .B(\B_not[9] ), .CI(\carry[9] ), .CO(\carry[10] ), 
        .S(DIFF[9]) );
  fa1a1 U2_8 ( .A(A[8]), .B(\B_not[8] ), .CI(\carry[8] ), .CO(\carry[9] ), .S(
        DIFF[8]) );
  fa1a1 U2_5 ( .A(A[5]), .B(\B_not[5] ), .CI(\carry[5] ), .CO(\carry[6] ), .S(
        DIFF[5]) );
  fa1a1 U2_4 ( .A(A[4]), .B(\B_not[4] ), .CI(\carry[4] ), .CO(\carry[5] ), .S(
        DIFF[4]) );
  fa1a1 U2_1 ( .A(A[1]), .B(\B_not[1] ), .CI(\carry[1] ), .CO(\carry[2] ), .S(
        DIFF[1]) );
  xor3a3 U2_29 ( .A(A[29]), .B(\B_not[29] ), .C(\carry[29] ), .Y(DIFF[29]) );
  or2a1 U1 ( .A(A[0]), .B(\B_not[0] ), .Y(\carry[1] ) );
  xor2a1 U2 ( .A(n1), .B(\B_not[0] ), .Y(DIFF[0]) );
  inv1a1 U3 ( .A(A[0]), .Y(n1) );
  inv1a1 U4 ( .A(B[9]), .Y(\B_not[9] ) );
  inv1a1 U5 ( .A(B[8]), .Y(\B_not[8] ) );
  inv1a1 U6 ( .A(B[7]), .Y(\B_not[7] ) );
  inv1a1 U7 ( .A(B[6]), .Y(\B_not[6] ) );
  inv1a1 U8 ( .A(B[5]), .Y(\B_not[5] ) );
  inv1a1 U9 ( .A(B[4]), .Y(\B_not[4] ) );
  inv1a1 U10 ( .A(B[3]), .Y(\B_not[3] ) );
  inv1a1 U11 ( .A(B[2]), .Y(\B_not[2] ) );
  inv1a1 U12 ( .A(B[29]), .Y(\B_not[29] ) );
  inv1a1 U13 ( .A(B[28]), .Y(\B_not[28] ) );
  inv1a1 U14 ( .A(B[27]), .Y(\B_not[27] ) );
  inv1a1 U15 ( .A(B[26]), .Y(\B_not[26] ) );
  inv1a1 U16 ( .A(B[25]), .Y(\B_not[25] ) );
  inv1a1 U17 ( .A(B[24]), .Y(\B_not[24] ) );
  inv1a1 U18 ( .A(B[23]), .Y(\B_not[23] ) );
  inv1a1 U19 ( .A(B[22]), .Y(\B_not[22] ) );
  inv1a1 U20 ( .A(B[21]), .Y(\B_not[21] ) );
  inv1a1 U21 ( .A(B[20]), .Y(\B_not[20] ) );
  inv1a1 U22 ( .A(B[1]), .Y(\B_not[1] ) );
  inv1a1 U23 ( .A(B[19]), .Y(\B_not[19] ) );
  inv1a1 U24 ( .A(B[18]), .Y(\B_not[18] ) );
  inv1a1 U25 ( .A(B[17]), .Y(\B_not[17] ) );
  inv1a1 U26 ( .A(B[16]), .Y(\B_not[16] ) );
  inv1a1 U27 ( .A(B[15]), .Y(\B_not[15] ) );
  inv1a1 U28 ( .A(B[14]), .Y(\B_not[14] ) );
  inv1a1 U29 ( .A(B[13]), .Y(\B_not[13] ) );
  inv1a1 U30 ( .A(B[12]), .Y(\B_not[12] ) );
  inv1a1 U31 ( .A(B[11]), .Y(\B_not[11] ) );
  inv1a1 U32 ( .A(B[10]), .Y(\B_not[10] ) );
  inv1a1 U33 ( .A(B[0]), .Y(\B_not[0] ) );
endmodule


module b14_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221;

  ao1f1 U1 ( .A(n1), .B(n2), .C(n3), .Y(LT) );
  oa1f1 U2 ( .A(n4), .B(n5), .C(n6), .Y(n2) );
  and2a3 U3 ( .A(B[30]), .B(n7), .Y(n6) );
  oa1f1 U4 ( .A(n8), .B(n9), .C(n10), .Y(n4) );
  oa1f1 U5 ( .A(n11), .B(n12), .C(n13), .Y(n8) );
  oa1f1 U6 ( .A(n14), .B(n15), .C(n16), .Y(n11) );
  inv1a1 U7 ( .A(n17), .Y(n16) );
  oa1f1 U8 ( .A(n18), .B(n19), .C(n20), .Y(n14) );
  oa1f1 U9 ( .A(n21), .B(n22), .C(n23), .Y(n18) );
  oa1f1 U10 ( .A(n24), .B(n25), .C(n26), .Y(n21) );
  oa1f1 U11 ( .A(n27), .B(n28), .C(n29), .Y(n24) );
  inv1a1 U12 ( .A(n30), .Y(n29) );
  oa1f1 U13 ( .A(n31), .B(n32), .C(n33), .Y(n27) );
  oa1f1 U14 ( .A(n34), .B(n35), .C(n36), .Y(n31) );
  oa1f1 U15 ( .A(n37), .B(n38), .C(n39), .Y(n34) );
  oa1f1 U16 ( .A(n40), .B(n41), .C(n42), .Y(n37) );
  inv1a1 U17 ( .A(n43), .Y(n42) );
  oa1f1 U18 ( .A(n44), .B(n45), .C(n46), .Y(n40) );
  oa1f1 U19 ( .A(n47), .B(n48), .C(n49), .Y(n44) );
  oa1f1 U20 ( .A(n50), .B(n51), .C(n52), .Y(n47) );
  oa1f1 U21 ( .A(n53), .B(n54), .C(n55), .Y(n50) );
  inv1a1 U22 ( .A(n56), .Y(n55) );
  oa1f1 U23 ( .A(n57), .B(n58), .C(n59), .Y(n53) );
  oa1f1 U24 ( .A(n60), .B(n61), .C(n62), .Y(n57) );
  oa1f1 U25 ( .A(n63), .B(n64), .C(n65), .Y(n60) );
  oa1f1 U26 ( .A(n66), .B(n67), .C(n68), .Y(n63) );
  inv1a1 U27 ( .A(n69), .Y(n68) );
  oa1f1 U28 ( .A(n70), .B(n71), .C(n72), .Y(n66) );
  oa1f1 U29 ( .A(n73), .B(n74), .C(n75), .Y(n70) );
  oa1f1 U30 ( .A(n76), .B(n77), .C(n78), .Y(n73) );
  oa1f1 U31 ( .A(n79), .B(n80), .C(n81), .Y(n76) );
  inv1a1 U32 ( .A(n82), .Y(n81) );
  oa1f1 U33 ( .A(n83), .B(n84), .C(n85), .Y(n79) );
  oa1f1 U34 ( .A(n86), .B(n87), .C(n88), .Y(n83) );
  oa1f1 U35 ( .A(n89), .B(n90), .C(n91), .Y(n86) );
  oa1f1 U36 ( .A(n92), .B(n93), .C(n94), .Y(n89) );
  inv1a1 U37 ( .A(n95), .Y(n94) );
  oa1f1 U38 ( .A(n96), .B(n97), .C(n98), .Y(n92) );
  oa1f1 U39 ( .A(A[1]), .B(n99), .C(n100), .Y(n96) );
  inv1a1 U40 ( .A(n101), .Y(n100) );
  ao1f1 U41 ( .A(n99), .B(A[1]), .C(n102), .Y(n101) );
  or2a1 U42 ( .A(A[0]), .B(n103), .Y(n99) );
  ao1a1 U43 ( .A(n104), .B(n3), .C(n1), .Y(GT) );
  and2a3 U44 ( .A(n105), .B(B[31]), .Y(n1) );
  or2a1 U45 ( .A(B[31]), .B(n105), .Y(n3) );
  inv1a1 U46 ( .A(A[31]), .Y(n105) );
  ao1f1 U47 ( .A(n106), .B(n107), .C(n108), .Y(n104) );
  or2a1 U48 ( .A(B[30]), .B(n7), .Y(n108) );
  ao1f1 U49 ( .A(n109), .B(n110), .C(n9), .Y(n107) );
  or2a1 U50 ( .A(A[29]), .B(n111), .Y(n9) );
  or2a1 U51 ( .A(n112), .B(n10), .Y(n110) );
  and2a3 U52 ( .A(n111), .B(A[29]), .Y(n10) );
  inv1a1 U53 ( .A(B[29]), .Y(n111) );
  and3a1 U54 ( .A(n113), .B(n15), .C(n12), .Y(n109) );
  inv1a1 U55 ( .A(n114), .Y(n12) );
  or2a1 U56 ( .A(n13), .B(n112), .Y(n114) );
  and2a3 U57 ( .A(n115), .B(A[28]), .Y(n112) );
  inv1a1 U58 ( .A(B[28]), .Y(n115) );
  and2a3 U59 ( .A(n116), .B(B[28]), .Y(n13) );
  inv1a1 U60 ( .A(A[28]), .Y(n116) );
  inv1a1 U61 ( .A(n117), .Y(n15) );
  and2a3 U62 ( .A(n118), .B(B[27]), .Y(n117) );
  ao1f1 U63 ( .A(n119), .B(n120), .C(n121), .Y(n113) );
  and2a3 U64 ( .A(n17), .B(n122), .Y(n121) );
  or2a1 U65 ( .A(B[27]), .B(n118), .Y(n17) );
  inv1a1 U66 ( .A(A[27]), .Y(n118) );
  ao1f1 U67 ( .A(n123), .B(n124), .C(n22), .Y(n120) );
  or2a1 U68 ( .A(A[25]), .B(n125), .Y(n22) );
  or2a1 U69 ( .A(n126), .B(n23), .Y(n124) );
  and2a3 U70 ( .A(n125), .B(A[25]), .Y(n23) );
  inv1a1 U71 ( .A(B[25]), .Y(n125) );
  and3a1 U72 ( .A(n127), .B(n28), .C(n25), .Y(n123) );
  inv1a1 U73 ( .A(n128), .Y(n25) );
  or2a1 U74 ( .A(n26), .B(n126), .Y(n128) );
  and2a3 U75 ( .A(n129), .B(A[24]), .Y(n126) );
  inv1a1 U76 ( .A(B[24]), .Y(n129) );
  and2a3 U77 ( .A(n130), .B(B[24]), .Y(n26) );
  inv1a1 U78 ( .A(A[24]), .Y(n130) );
  inv1a1 U79 ( .A(n131), .Y(n28) );
  and2a3 U80 ( .A(n132), .B(B[23]), .Y(n131) );
  ao1f1 U81 ( .A(n133), .B(n134), .C(n135), .Y(n127) );
  and2a3 U82 ( .A(n30), .B(n136), .Y(n135) );
  or2a1 U83 ( .A(B[23]), .B(n132), .Y(n30) );
  inv1a1 U84 ( .A(A[23]), .Y(n132) );
  ao1f1 U85 ( .A(n137), .B(n138), .C(n35), .Y(n134) );
  or2a1 U86 ( .A(A[21]), .B(n139), .Y(n35) );
  or2a1 U87 ( .A(n140), .B(n36), .Y(n138) );
  and2a3 U88 ( .A(n139), .B(A[21]), .Y(n36) );
  inv1a1 U89 ( .A(B[21]), .Y(n139) );
  and3a1 U90 ( .A(n141), .B(n41), .C(n38), .Y(n137) );
  inv1a1 U91 ( .A(n142), .Y(n38) );
  or2a1 U92 ( .A(n39), .B(n140), .Y(n142) );
  and2a3 U93 ( .A(n143), .B(A[20]), .Y(n140) );
  inv1a1 U94 ( .A(B[20]), .Y(n143) );
  and2a3 U95 ( .A(n144), .B(B[20]), .Y(n39) );
  inv1a1 U96 ( .A(A[20]), .Y(n144) );
  inv1a1 U97 ( .A(n145), .Y(n41) );
  and2a3 U98 ( .A(n146), .B(B[19]), .Y(n145) );
  ao1f1 U99 ( .A(n147), .B(n148), .C(n149), .Y(n141) );
  and2a3 U100 ( .A(n43), .B(n150), .Y(n149) );
  or2a1 U101 ( .A(B[19]), .B(n146), .Y(n43) );
  inv1a1 U102 ( .A(A[19]), .Y(n146) );
  ao1f1 U103 ( .A(n151), .B(n152), .C(n48), .Y(n148) );
  or2a1 U104 ( .A(A[17]), .B(n153), .Y(n48) );
  or2a1 U105 ( .A(n154), .B(n49), .Y(n152) );
  and2a3 U106 ( .A(n153), .B(A[17]), .Y(n49) );
  inv1a1 U107 ( .A(B[17]), .Y(n153) );
  and3a1 U108 ( .A(n155), .B(n54), .C(n51), .Y(n151) );
  inv1a1 U109 ( .A(n156), .Y(n51) );
  or2a1 U110 ( .A(n52), .B(n154), .Y(n156) );
  and2a3 U111 ( .A(n157), .B(A[16]), .Y(n154) );
  inv1a1 U112 ( .A(B[16]), .Y(n157) );
  and2a3 U113 ( .A(n158), .B(B[16]), .Y(n52) );
  inv1a1 U114 ( .A(A[16]), .Y(n158) );
  inv1a1 U115 ( .A(n159), .Y(n54) );
  and2a3 U116 ( .A(n160), .B(B[15]), .Y(n159) );
  ao1f1 U117 ( .A(n161), .B(n162), .C(n163), .Y(n155) );
  and2a3 U118 ( .A(n56), .B(n164), .Y(n163) );
  or2a1 U119 ( .A(B[15]), .B(n160), .Y(n56) );
  inv1a1 U120 ( .A(A[15]), .Y(n160) );
  ao1f1 U121 ( .A(n165), .B(n166), .C(n61), .Y(n162) );
  or2a1 U122 ( .A(A[13]), .B(n167), .Y(n61) );
  or2a1 U123 ( .A(n168), .B(n62), .Y(n166) );
  and2a3 U124 ( .A(n167), .B(A[13]), .Y(n62) );
  inv1a1 U125 ( .A(B[13]), .Y(n167) );
  and3a1 U126 ( .A(n169), .B(n67), .C(n64), .Y(n165) );
  inv1a1 U127 ( .A(n170), .Y(n64) );
  or2a1 U128 ( .A(n65), .B(n168), .Y(n170) );
  and2a3 U129 ( .A(n171), .B(A[12]), .Y(n168) );
  inv1a1 U130 ( .A(B[12]), .Y(n171) );
  and2a3 U131 ( .A(n172), .B(B[12]), .Y(n65) );
  inv1a1 U132 ( .A(A[12]), .Y(n172) );
  inv1a1 U133 ( .A(n173), .Y(n67) );
  and2a3 U134 ( .A(n174), .B(B[11]), .Y(n173) );
  ao1f1 U135 ( .A(n175), .B(n176), .C(n177), .Y(n169) );
  and2a3 U136 ( .A(n69), .B(n178), .Y(n177) );
  or2a1 U137 ( .A(B[11]), .B(n174), .Y(n69) );
  inv1a1 U138 ( .A(A[11]), .Y(n174) );
  ao1f1 U139 ( .A(n179), .B(n180), .C(n74), .Y(n176) );
  or2a1 U140 ( .A(A[9]), .B(n181), .Y(n74) );
  or2a1 U141 ( .A(n182), .B(n75), .Y(n180) );
  and2a3 U142 ( .A(n181), .B(A[9]), .Y(n75) );
  inv1a1 U143 ( .A(B[9]), .Y(n181) );
  and3a1 U144 ( .A(n183), .B(n80), .C(n77), .Y(n179) );
  inv1a1 U145 ( .A(n184), .Y(n77) );
  or2a1 U146 ( .A(n78), .B(n182), .Y(n184) );
  and2a3 U147 ( .A(n185), .B(A[8]), .Y(n182) );
  inv1a1 U148 ( .A(B[8]), .Y(n185) );
  and2a3 U149 ( .A(n186), .B(B[8]), .Y(n78) );
  inv1a1 U150 ( .A(A[8]), .Y(n186) );
  inv1a1 U151 ( .A(n187), .Y(n80) );
  and2a3 U152 ( .A(n188), .B(B[7]), .Y(n187) );
  ao1f1 U153 ( .A(n189), .B(n190), .C(n191), .Y(n183) );
  and2a3 U154 ( .A(n82), .B(n192), .Y(n191) );
  or2a1 U155 ( .A(B[7]), .B(n188), .Y(n82) );
  inv1a1 U156 ( .A(A[7]), .Y(n188) );
  ao1f1 U157 ( .A(n193), .B(n194), .C(n87), .Y(n190) );
  or2a1 U158 ( .A(A[5]), .B(n195), .Y(n87) );
  or2a1 U159 ( .A(n196), .B(n88), .Y(n194) );
  and2a3 U160 ( .A(n195), .B(A[5]), .Y(n88) );
  inv1a1 U161 ( .A(B[5]), .Y(n195) );
  and3a1 U162 ( .A(n197), .B(n93), .C(n90), .Y(n193) );
  inv1a1 U163 ( .A(n198), .Y(n90) );
  or2a1 U164 ( .A(n91), .B(n196), .Y(n198) );
  and2a3 U165 ( .A(n199), .B(A[4]), .Y(n196) );
  inv1a1 U166 ( .A(B[4]), .Y(n199) );
  and2a3 U167 ( .A(n200), .B(B[4]), .Y(n91) );
  inv1a1 U168 ( .A(A[4]), .Y(n200) );
  inv1a1 U169 ( .A(n201), .Y(n93) );
  and2a3 U170 ( .A(n202), .B(B[3]), .Y(n201) );
  ao1f1 U171 ( .A(n203), .B(n204), .C(n205), .Y(n197) );
  and2a3 U172 ( .A(n95), .B(n206), .Y(n205) );
  or2a1 U173 ( .A(B[3]), .B(n202), .Y(n95) );
  inv1a1 U174 ( .A(A[3]), .Y(n202) );
  fac2a1 U175 ( .A(A[1]), .B(n102), .CI(n207), .CO(n204) );
  and2a3 U176 ( .A(A[0]), .B(n103), .Y(n207) );
  inv1a1 U177 ( .A(B[0]), .Y(n103) );
  inv1a1 U178 ( .A(B[1]), .Y(n102) );
  inv1a1 U179 ( .A(n97), .Y(n203) );
  and2a3 U180 ( .A(n208), .B(n206), .Y(n97) );
  or2a1 U181 ( .A(B[2]), .B(n209), .Y(n206) );
  inv1a1 U182 ( .A(n98), .Y(n208) );
  and2a3 U183 ( .A(n209), .B(B[2]), .Y(n98) );
  inv1a1 U184 ( .A(A[2]), .Y(n209) );
  inv1a1 U185 ( .A(n84), .Y(n189) );
  and2a3 U186 ( .A(n210), .B(n192), .Y(n84) );
  or2a1 U187 ( .A(B[6]), .B(n211), .Y(n192) );
  inv1a1 U188 ( .A(n85), .Y(n210) );
  and2a3 U189 ( .A(n211), .B(B[6]), .Y(n85) );
  inv1a1 U190 ( .A(A[6]), .Y(n211) );
  inv1a1 U191 ( .A(n71), .Y(n175) );
  and2a3 U192 ( .A(n212), .B(n178), .Y(n71) );
  or2a1 U193 ( .A(B[10]), .B(n213), .Y(n178) );
  inv1a1 U194 ( .A(n72), .Y(n212) );
  and2a3 U195 ( .A(n213), .B(B[10]), .Y(n72) );
  inv1a1 U196 ( .A(A[10]), .Y(n213) );
  inv1a1 U197 ( .A(n58), .Y(n161) );
  and2a3 U198 ( .A(n214), .B(n164), .Y(n58) );
  or2a1 U199 ( .A(B[14]), .B(n215), .Y(n164) );
  inv1a1 U200 ( .A(n59), .Y(n214) );
  and2a3 U201 ( .A(n215), .B(B[14]), .Y(n59) );
  inv1a1 U202 ( .A(A[14]), .Y(n215) );
  inv1a1 U203 ( .A(n45), .Y(n147) );
  and2a3 U204 ( .A(n216), .B(n150), .Y(n45) );
  or2a1 U205 ( .A(B[18]), .B(n217), .Y(n150) );
  inv1a1 U206 ( .A(n46), .Y(n216) );
  and2a3 U207 ( .A(n217), .B(B[18]), .Y(n46) );
  inv1a1 U208 ( .A(A[18]), .Y(n217) );
  inv1a1 U209 ( .A(n32), .Y(n133) );
  and2a3 U210 ( .A(n218), .B(n136), .Y(n32) );
  or2a1 U211 ( .A(B[22]), .B(n219), .Y(n136) );
  inv1a1 U212 ( .A(n33), .Y(n218) );
  and2a3 U213 ( .A(n219), .B(B[22]), .Y(n33) );
  inv1a1 U214 ( .A(A[22]), .Y(n219) );
  inv1a1 U215 ( .A(n19), .Y(n119) );
  and2a3 U216 ( .A(n220), .B(n122), .Y(n19) );
  or2a1 U217 ( .A(B[26]), .B(n221), .Y(n122) );
  inv1a1 U218 ( .A(n20), .Y(n220) );
  and2a3 U219 ( .A(n221), .B(B[26]), .Y(n20) );
  inv1a1 U220 ( .A(A[26]), .Y(n221) );
  inv1a1 U221 ( .A(n5), .Y(n106) );
  xor2a1 U222 ( .A(n7), .B(B[30]), .Y(n5) );
  inv1a1 U223 ( .A(A[30]), .Y(n7) );
endmodule


module b14_DW01_addsub_2 ( A, B, CI, ADD_SUB, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ,
         \carry[1] , \carry[0] , \B_AS[31] , \B_AS[30] , \B_AS[18] ,
         \B_AS[17] , \B_AS[16] , \B_AS[15] , \B_AS[14] , \B_AS[13] ,
         \B_AS[12] , \B_AS[11] , \B_AS[10] , \B_AS[9] , \B_AS[8] , \B_AS[7] ,
         \B_AS[6] , \B_AS[5] , \B_AS[4] , \B_AS[3] , \B_AS[2] , \B_AS[1] ,
         \B_AS[0] ;
  assign \carry[0]  = ADD_SUB;

  fa1a1 U1_1 ( .A(A[1]), .B(\B_AS[1] ), .CI(\carry[1] ), .CO(\carry[2] ), .S(
        SUM[1]) );
  fa1a1 U1_2 ( .A(A[2]), .B(\B_AS[2] ), .CI(\carry[2] ), .CO(\carry[3] ), .S(
        SUM[2]) );
  fa1a1 U1_3 ( .A(A[3]), .B(\B_AS[3] ), .CI(\carry[3] ), .CO(\carry[4] ), .S(
        SUM[3]) );
  fa1a1 U1_4 ( .A(A[4]), .B(\B_AS[4] ), .CI(\carry[4] ), .CO(\carry[5] ), .S(
        SUM[4]) );
  fa1a1 U1_5 ( .A(A[5]), .B(\B_AS[5] ), .CI(\carry[5] ), .CO(\carry[6] ), .S(
        SUM[5]) );
  fa1a1 U1_6 ( .A(A[6]), .B(\B_AS[6] ), .CI(\carry[6] ), .CO(\carry[7] ), .S(
        SUM[6]) );
  fa1a1 U1_7 ( .A(A[7]), .B(\B_AS[7] ), .CI(\carry[7] ), .CO(\carry[8] ), .S(
        SUM[7]) );
  fa1a1 U1_8 ( .A(A[8]), .B(\B_AS[8] ), .CI(\carry[8] ), .CO(\carry[9] ), .S(
        SUM[8]) );
  fa1a1 U1_9 ( .A(A[9]), .B(\B_AS[9] ), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  fa1a1 U1_10 ( .A(A[10]), .B(\B_AS[10] ), .CI(\carry[10] ), .CO(\carry[11] ), 
        .S(SUM[10]) );
  fa1a1 U1_11 ( .A(A[11]), .B(\B_AS[11] ), .CI(\carry[11] ), .CO(\carry[12] ), 
        .S(SUM[11]) );
  fa1a1 U1_12 ( .A(A[12]), .B(\B_AS[12] ), .CI(\carry[12] ), .CO(\carry[13] ), 
        .S(SUM[12]) );
  fa1a1 U1_13 ( .A(A[13]), .B(\B_AS[13] ), .CI(\carry[13] ), .CO(\carry[14] ), 
        .S(SUM[13]) );
  fa1a1 U1_14 ( .A(A[14]), .B(\B_AS[14] ), .CI(\carry[14] ), .CO(\carry[15] ), 
        .S(SUM[14]) );
  fa1a1 U1_15 ( .A(A[15]), .B(\B_AS[15] ), .CI(\carry[15] ), .CO(\carry[16] ), 
        .S(SUM[15]) );
  fa1a1 U1_16 ( .A(A[16]), .B(\B_AS[16] ), .CI(\carry[16] ), .CO(\carry[17] ), 
        .S(SUM[16]) );
  fa1a1 U1_17 ( .A(A[17]), .B(\B_AS[17] ), .CI(\carry[17] ), .CO(\carry[18] ), 
        .S(SUM[17]) );
  fa1a1 U1_18 ( .A(A[18]), .B(\B_AS[18] ), .CI(\carry[18] ), .CO(\carry[19] ), 
        .S(SUM[18]) );
  fa1a1 U1_30 ( .A(A[30]), .B(\B_AS[30] ), .CI(\carry[30] ), .CO(\carry[31] ), 
        .S(SUM[30]) );
  fa1a1 U1_0 ( .A(A[0]), .B(\B_AS[0] ), .CI(\carry[0] ), .CO(\carry[1] ), .S(
        SUM[0]) );
  fa1a1 U1_28 ( .A(A[28]), .B(\B_AS[31] ), .CI(\carry[28] ), .CO(\carry[29] ), 
        .S(SUM[28]) );
  fa1a1 U1_19 ( .A(A[19]), .B(\B_AS[31] ), .CI(\carry[19] ), .CO(\carry[20] ), 
        .S(SUM[19]) );
  fa1a1 U1_20 ( .A(A[20]), .B(\B_AS[31] ), .CI(\carry[20] ), .CO(\carry[21] ), 
        .S(SUM[20]) );
  fa1a1 U1_21 ( .A(A[21]), .B(\B_AS[31] ), .CI(\carry[21] ), .CO(\carry[22] ), 
        .S(SUM[21]) );
  fa1a1 U1_22 ( .A(A[22]), .B(\B_AS[31] ), .CI(\carry[22] ), .CO(\carry[23] ), 
        .S(SUM[22]) );
  fa1a1 U1_23 ( .A(A[23]), .B(\B_AS[31] ), .CI(\carry[23] ), .CO(\carry[24] ), 
        .S(SUM[23]) );
  fa1a1 U1_24 ( .A(A[24]), .B(\B_AS[31] ), .CI(\carry[24] ), .CO(\carry[25] ), 
        .S(SUM[24]) );
  fa1a1 U1_25 ( .A(A[25]), .B(\B_AS[31] ), .CI(\carry[25] ), .CO(\carry[26] ), 
        .S(SUM[25]) );
  fa1a1 U1_26 ( .A(A[26]), .B(\B_AS[31] ), .CI(\carry[26] ), .CO(\carry[27] ), 
        .S(SUM[26]) );
  fa1a1 U1_27 ( .A(A[27]), .B(\B_AS[31] ), .CI(\carry[27] ), .CO(\carry[28] ), 
        .S(SUM[27]) );
  fa1a1 U1_29 ( .A(A[29]), .B(\B_AS[31] ), .CI(\carry[29] ), .CO(\carry[30] ), 
        .S(SUM[29]) );
  xor3a3 U1_31 ( .A(A[31]), .B(\B_AS[31] ), .C(\carry[31] ), .Y(SUM[31]) );
  xor2a6 U1 ( .A(\carry[0] ), .B(B[31]), .Y(\B_AS[31] ) );
  xor2a1 U2 ( .A(B[9]), .B(\carry[0] ), .Y(\B_AS[9] ) );
  xor2a1 U3 ( .A(B[8]), .B(\carry[0] ), .Y(\B_AS[8] ) );
  xor2a1 U4 ( .A(B[7]), .B(\carry[0] ), .Y(\B_AS[7] ) );
  xor2a1 U5 ( .A(B[6]), .B(\carry[0] ), .Y(\B_AS[6] ) );
  xor2a1 U6 ( .A(B[5]), .B(\carry[0] ), .Y(\B_AS[5] ) );
  xor2a1 U7 ( .A(B[4]), .B(\carry[0] ), .Y(\B_AS[4] ) );
  xor2a1 U8 ( .A(B[3]), .B(\carry[0] ), .Y(\B_AS[3] ) );
  xor2a1 U9 ( .A(B[30]), .B(\carry[0] ), .Y(\B_AS[30] ) );
  xor2a1 U10 ( .A(B[2]), .B(\carry[0] ), .Y(\B_AS[2] ) );
  xor2a1 U11 ( .A(B[1]), .B(\carry[0] ), .Y(\B_AS[1] ) );
  xor2a1 U12 ( .A(B[18]), .B(\carry[0] ), .Y(\B_AS[18] ) );
  xor2a1 U13 ( .A(B[17]), .B(\carry[0] ), .Y(\B_AS[17] ) );
  xor2a1 U14 ( .A(B[16]), .B(\carry[0] ), .Y(\B_AS[16] ) );
  xor2a1 U15 ( .A(B[15]), .B(\carry[0] ), .Y(\B_AS[15] ) );
  xor2a1 U16 ( .A(B[14]), .B(\carry[0] ), .Y(\B_AS[14] ) );
  xor2a1 U17 ( .A(B[13]), .B(\carry[0] ), .Y(\B_AS[13] ) );
  xor2a1 U18 ( .A(B[12]), .B(\carry[0] ), .Y(\B_AS[12] ) );
  xor2a1 U19 ( .A(B[11]), .B(\carry[0] ), .Y(\B_AS[11] ) );
  xor2a1 U20 ( .A(B[10]), .B(\carry[0] ), .Y(\B_AS[10] ) );
  xor2a1 U21 ( .A(B[0]), .B(\carry[0] ), .Y(\B_AS[0] ) );
endmodule


module b14_DW01_cmp2_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [31:0] A;
  input [31:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;

  ao1f1 U1 ( .A(n1), .B(n2), .C(n3), .Y(LT_LE) );
  or2a1 U2 ( .A(B[31]), .B(n4), .Y(n3) );
  oa1f1 U3 ( .A(n5), .B(n6), .C(n7), .Y(n2) );
  and2a3 U4 ( .A(B[30]), .B(n8), .Y(n7) );
  or2a1 U5 ( .A(B[30]), .B(n8), .Y(n6) );
  inv1a1 U6 ( .A(A[30]), .Y(n8) );
  oa1f1 U7 ( .A(n9), .B(n10), .C(n11), .Y(n5) );
  and2a3 U8 ( .A(A[29]), .B(n12), .Y(n11) );
  or2a1 U9 ( .A(A[29]), .B(n12), .Y(n10) );
  inv1a1 U10 ( .A(B[29]), .Y(n12) );
  oa1f1 U11 ( .A(n13), .B(n14), .C(n15), .Y(n9) );
  and2a3 U12 ( .A(B[28]), .B(n16), .Y(n15) );
  or2a1 U13 ( .A(B[28]), .B(n16), .Y(n14) );
  inv1a1 U14 ( .A(A[28]), .Y(n16) );
  oa1f1 U15 ( .A(n17), .B(n18), .C(n19), .Y(n13) );
  and2a3 U16 ( .A(A[27]), .B(n20), .Y(n19) );
  or2a1 U17 ( .A(A[27]), .B(n20), .Y(n18) );
  inv1a1 U18 ( .A(B[27]), .Y(n20) );
  oa1f1 U19 ( .A(n21), .B(n22), .C(n23), .Y(n17) );
  and2a3 U20 ( .A(B[26]), .B(n24), .Y(n23) );
  or2a1 U21 ( .A(B[26]), .B(n24), .Y(n22) );
  inv1a1 U22 ( .A(A[26]), .Y(n24) );
  oa1f1 U23 ( .A(n25), .B(n26), .C(n27), .Y(n21) );
  and2a3 U24 ( .A(A[25]), .B(n28), .Y(n27) );
  or2a1 U25 ( .A(A[25]), .B(n28), .Y(n26) );
  inv1a1 U26 ( .A(B[25]), .Y(n28) );
  oa1f1 U27 ( .A(n29), .B(n30), .C(n31), .Y(n25) );
  and2a3 U28 ( .A(B[24]), .B(n32), .Y(n31) );
  or2a1 U29 ( .A(B[24]), .B(n32), .Y(n30) );
  inv1a1 U30 ( .A(A[24]), .Y(n32) );
  oa1f1 U31 ( .A(n33), .B(n34), .C(n35), .Y(n29) );
  and2a3 U32 ( .A(A[23]), .B(n36), .Y(n35) );
  or2a1 U33 ( .A(A[23]), .B(n36), .Y(n34) );
  inv1a1 U34 ( .A(B[23]), .Y(n36) );
  oa1f1 U35 ( .A(n37), .B(n38), .C(n39), .Y(n33) );
  and2a3 U36 ( .A(B[22]), .B(n40), .Y(n39) );
  or2a1 U37 ( .A(B[22]), .B(n40), .Y(n38) );
  inv1a1 U38 ( .A(A[22]), .Y(n40) );
  oa1f1 U39 ( .A(n41), .B(n42), .C(n43), .Y(n37) );
  and2a3 U40 ( .A(A[21]), .B(n44), .Y(n43) );
  or2a1 U41 ( .A(A[21]), .B(n44), .Y(n42) );
  inv1a1 U42 ( .A(B[21]), .Y(n44) );
  oa1f1 U43 ( .A(n45), .B(n46), .C(n47), .Y(n41) );
  and2a3 U44 ( .A(B[20]), .B(n48), .Y(n47) );
  or2a1 U45 ( .A(B[20]), .B(n48), .Y(n46) );
  inv1a1 U46 ( .A(A[20]), .Y(n48) );
  oa1f1 U47 ( .A(n49), .B(n50), .C(n51), .Y(n45) );
  and2a3 U48 ( .A(A[19]), .B(n52), .Y(n51) );
  or2a1 U49 ( .A(A[19]), .B(n52), .Y(n50) );
  inv1a1 U50 ( .A(B[19]), .Y(n52) );
  oa1f1 U51 ( .A(n53), .B(n54), .C(n55), .Y(n49) );
  and2a3 U52 ( .A(B[18]), .B(n56), .Y(n55) );
  or2a1 U53 ( .A(B[18]), .B(n56), .Y(n54) );
  inv1a1 U54 ( .A(A[18]), .Y(n56) );
  oa1f1 U55 ( .A(n57), .B(n58), .C(n59), .Y(n53) );
  and2a3 U56 ( .A(A[17]), .B(n60), .Y(n59) );
  or2a1 U57 ( .A(A[17]), .B(n60), .Y(n58) );
  inv1a1 U58 ( .A(B[17]), .Y(n60) );
  oa1f1 U59 ( .A(n61), .B(n62), .C(n63), .Y(n57) );
  and2a3 U60 ( .A(B[16]), .B(n64), .Y(n63) );
  or2a1 U61 ( .A(B[16]), .B(n64), .Y(n62) );
  inv1a1 U62 ( .A(A[16]), .Y(n64) );
  oa1f1 U63 ( .A(n65), .B(n66), .C(n67), .Y(n61) );
  and2a3 U64 ( .A(A[15]), .B(n68), .Y(n67) );
  or2a1 U65 ( .A(A[15]), .B(n68), .Y(n66) );
  inv1a1 U66 ( .A(B[15]), .Y(n68) );
  oa1f1 U67 ( .A(n69), .B(n70), .C(n71), .Y(n65) );
  and2a3 U68 ( .A(B[14]), .B(n72), .Y(n71) );
  or2a1 U69 ( .A(B[14]), .B(n72), .Y(n70) );
  inv1a1 U70 ( .A(A[14]), .Y(n72) );
  oa1f1 U71 ( .A(n73), .B(n74), .C(n75), .Y(n69) );
  and2a3 U72 ( .A(A[13]), .B(n76), .Y(n75) );
  or2a1 U73 ( .A(A[13]), .B(n76), .Y(n74) );
  inv1a1 U74 ( .A(B[13]), .Y(n76) );
  oa1f1 U75 ( .A(n77), .B(n78), .C(n79), .Y(n73) );
  and2a3 U76 ( .A(B[12]), .B(n80), .Y(n79) );
  or2a1 U77 ( .A(B[12]), .B(n80), .Y(n78) );
  inv1a1 U78 ( .A(A[12]), .Y(n80) );
  oa1f1 U79 ( .A(n81), .B(n82), .C(n83), .Y(n77) );
  and2a3 U80 ( .A(A[11]), .B(n84), .Y(n83) );
  or2a1 U81 ( .A(A[11]), .B(n84), .Y(n82) );
  inv1a1 U82 ( .A(B[11]), .Y(n84) );
  oa1f1 U83 ( .A(n85), .B(n86), .C(n87), .Y(n81) );
  and2a3 U84 ( .A(B[10]), .B(n88), .Y(n87) );
  inv1a1 U85 ( .A(A[10]), .Y(n88) );
  or2a1 U86 ( .A(B[9]), .B(n89), .Y(n86) );
  oa1f1 U87 ( .A(n90), .B(n91), .C(n92), .Y(n85) );
  and2a3 U88 ( .A(A[10]), .B(n93), .Y(n92) );
  inv1a1 U89 ( .A(B[10]), .Y(n93) );
  inv1a1 U90 ( .A(n94), .Y(n91) );
  and2a3 U91 ( .A(n89), .B(B[9]), .Y(n94) );
  inv1a1 U92 ( .A(A[9]), .Y(n89) );
  oa1f1 U93 ( .A(n95), .B(n96), .C(n97), .Y(n90) );
  and2a3 U94 ( .A(B[8]), .B(n98), .Y(n97) );
  or2a1 U95 ( .A(B[8]), .B(n98), .Y(n96) );
  inv1a1 U96 ( .A(A[8]), .Y(n98) );
  oa1f1 U97 ( .A(n99), .B(n100), .C(n101), .Y(n95) );
  and2a3 U98 ( .A(A[7]), .B(n102), .Y(n101) );
  or2a1 U99 ( .A(A[7]), .B(n102), .Y(n100) );
  inv1a1 U100 ( .A(B[7]), .Y(n102) );
  oa1f1 U101 ( .A(n103), .B(n104), .C(n105), .Y(n99) );
  and2a3 U102 ( .A(B[6]), .B(n106), .Y(n105) );
  or2a1 U103 ( .A(B[6]), .B(n106), .Y(n104) );
  inv1a1 U104 ( .A(A[6]), .Y(n106) );
  oa1f1 U105 ( .A(n107), .B(n108), .C(n109), .Y(n103) );
  and2a3 U106 ( .A(A[5]), .B(n110), .Y(n109) );
  or2a1 U107 ( .A(A[5]), .B(n110), .Y(n108) );
  inv1a1 U108 ( .A(B[5]), .Y(n110) );
  oa1f1 U109 ( .A(n111), .B(n112), .C(n113), .Y(n107) );
  and2a3 U110 ( .A(B[4]), .B(n114), .Y(n113) );
  or2a1 U111 ( .A(B[4]), .B(n114), .Y(n112) );
  inv1a1 U112 ( .A(A[4]), .Y(n114) );
  oa1f1 U113 ( .A(n115), .B(n116), .C(n117), .Y(n111) );
  and2a3 U114 ( .A(A[3]), .B(n118), .Y(n117) );
  or2a1 U115 ( .A(A[3]), .B(n118), .Y(n116) );
  inv1a1 U116 ( .A(B[3]), .Y(n118) );
  oa1f1 U117 ( .A(n119), .B(n120), .C(n121), .Y(n115) );
  and2a3 U118 ( .A(B[2]), .B(n122), .Y(n121) );
  or2a1 U119 ( .A(B[2]), .B(n122), .Y(n120) );
  inv1a1 U120 ( .A(A[2]), .Y(n122) );
  oa1f1 U121 ( .A(A[1]), .B(n123), .C(n124), .Y(n119) );
  oa1f1 U122 ( .A(n125), .B(n126), .C(B[1]), .Y(n124) );
  inv1a1 U123 ( .A(A[1]), .Y(n126) );
  inv1a1 U124 ( .A(n125), .Y(n123) );
  and2a3 U125 ( .A(n127), .B(B[0]), .Y(n125) );
  inv1a1 U126 ( .A(A[0]), .Y(n127) );
  and2a3 U127 ( .A(B[31]), .B(n4), .Y(n1) );
  inv1a1 U128 ( .A(A[31]), .Y(n4) );
endmodule


module b14_DW01_addsub_1 ( A, B, CI, ADD_SUB, SUM, CO );
  input [28:0] A;
  input [28:0] B;
  output [28:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   \carry[28] , \carry[27] , \carry[26] , \carry[25] , \carry[24] ,
         \carry[23] , \carry[22] , \carry[21] , \carry[20] , \carry[19] ,
         \carry[18] , \carry[17] , \carry[16] , \carry[15] , \carry[14] ,
         \carry[13] , \carry[12] , \carry[11] , \carry[10] , \carry[9] ,
         \carry[8] , \carry[7] , \carry[6] , \carry[5] , \carry[4] ,
         \carry[3] , \carry[2] , \carry[1] , \carry[0] , \B_AS[28] ,
         \B_AS[27] , \B_AS[26] , \B_AS[25] , \B_AS[24] , \B_AS[23] ,
         \B_AS[22] , \B_AS[21] , \B_AS[20] , \B_AS[19] , \B_AS[18] ,
         \B_AS[17] , \B_AS[16] , \B_AS[15] , \B_AS[14] , \B_AS[13] ,
         \B_AS[12] , \B_AS[11] , \B_AS[10] , \B_AS[9] , \B_AS[8] , \B_AS[7] ,
         \B_AS[6] , \B_AS[5] , \B_AS[4] , \B_AS[3] , \B_AS[2] , \B_AS[1] ,
         \B_AS[0] ;
  assign \carry[0]  = ADD_SUB;

  xor3a3 U1_28 ( .A(A[28]), .B(\B_AS[28] ), .C(\carry[28] ), .Y(SUM[28]) );
  fa1a1 U1_1 ( .A(A[1]), .B(\B_AS[1] ), .CI(\carry[1] ), .CO(\carry[2] ), .S(
        SUM[1]) );
  fa1a1 U1_2 ( .A(A[2]), .B(\B_AS[2] ), .CI(\carry[2] ), .CO(\carry[3] ), .S(
        SUM[2]) );
  fa1a1 U1_3 ( .A(A[3]), .B(\B_AS[3] ), .CI(\carry[3] ), .CO(\carry[4] ), .S(
        SUM[3]) );
  fa1a1 U1_4 ( .A(A[4]), .B(\B_AS[4] ), .CI(\carry[4] ), .CO(\carry[5] ), .S(
        SUM[4]) );
  fa1a1 U1_5 ( .A(A[5]), .B(\B_AS[5] ), .CI(\carry[5] ), .CO(\carry[6] ), .S(
        SUM[5]) );
  fa1a1 U1_6 ( .A(A[6]), .B(\B_AS[6] ), .CI(\carry[6] ), .CO(\carry[7] ), .S(
        SUM[6]) );
  fa1a1 U1_7 ( .A(A[7]), .B(\B_AS[7] ), .CI(\carry[7] ), .CO(\carry[8] ), .S(
        SUM[7]) );
  fa1a1 U1_8 ( .A(A[8]), .B(\B_AS[8] ), .CI(\carry[8] ), .CO(\carry[9] ), .S(
        SUM[8]) );
  fa1a1 U1_9 ( .A(A[9]), .B(\B_AS[9] ), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  fa1a1 U1_10 ( .A(A[10]), .B(\B_AS[10] ), .CI(\carry[10] ), .CO(\carry[11] ), 
        .S(SUM[10]) );
  fa1a1 U1_11 ( .A(A[11]), .B(\B_AS[11] ), .CI(\carry[11] ), .CO(\carry[12] ), 
        .S(SUM[11]) );
  fa1a1 U1_12 ( .A(A[12]), .B(\B_AS[12] ), .CI(\carry[12] ), .CO(\carry[13] ), 
        .S(SUM[12]) );
  fa1a1 U1_13 ( .A(A[13]), .B(\B_AS[13] ), .CI(\carry[13] ), .CO(\carry[14] ), 
        .S(SUM[13]) );
  fa1a1 U1_14 ( .A(A[14]), .B(\B_AS[14] ), .CI(\carry[14] ), .CO(\carry[15] ), 
        .S(SUM[14]) );
  fa1a1 U1_15 ( .A(A[15]), .B(\B_AS[15] ), .CI(\carry[15] ), .CO(\carry[16] ), 
        .S(SUM[15]) );
  fa1a1 U1_16 ( .A(A[16]), .B(\B_AS[16] ), .CI(\carry[16] ), .CO(\carry[17] ), 
        .S(SUM[16]) );
  fa1a1 U1_17 ( .A(A[17]), .B(\B_AS[17] ), .CI(\carry[17] ), .CO(\carry[18] ), 
        .S(SUM[17]) );
  fa1a1 U1_18 ( .A(A[18]), .B(\B_AS[18] ), .CI(\carry[18] ), .CO(\carry[19] ), 
        .S(SUM[18]) );
  fa1a1 U1_19 ( .A(A[19]), .B(\B_AS[19] ), .CI(\carry[19] ), .CO(\carry[20] ), 
        .S(SUM[19]) );
  fa1a1 U1_20 ( .A(A[20]), .B(\B_AS[20] ), .CI(\carry[20] ), .CO(\carry[21] ), 
        .S(SUM[20]) );
  fa1a1 U1_21 ( .A(A[21]), .B(\B_AS[21] ), .CI(\carry[21] ), .CO(\carry[22] ), 
        .S(SUM[21]) );
  fa1a1 U1_22 ( .A(A[22]), .B(\B_AS[22] ), .CI(\carry[22] ), .CO(\carry[23] ), 
        .S(SUM[22]) );
  fa1a1 U1_23 ( .A(A[23]), .B(\B_AS[23] ), .CI(\carry[23] ), .CO(\carry[24] ), 
        .S(SUM[23]) );
  fa1a1 U1_24 ( .A(A[24]), .B(\B_AS[24] ), .CI(\carry[24] ), .CO(\carry[25] ), 
        .S(SUM[24]) );
  fa1a1 U1_25 ( .A(A[25]), .B(\B_AS[25] ), .CI(\carry[25] ), .CO(\carry[26] ), 
        .S(SUM[25]) );
  fa1a1 U1_26 ( .A(A[26]), .B(\B_AS[26] ), .CI(\carry[26] ), .CO(\carry[27] ), 
        .S(SUM[26]) );
  fa1a1 U1_27 ( .A(A[27]), .B(\B_AS[27] ), .CI(\carry[27] ), .CO(\carry[28] ), 
        .S(SUM[27]) );
  fa1a1 U1_0 ( .A(A[0]), .B(\B_AS[0] ), .CI(\carry[0] ), .CO(\carry[1] ), .S(
        SUM[0]) );
  xor2a1 U1 ( .A(B[9]), .B(\carry[0] ), .Y(\B_AS[9] ) );
  xor2a1 U2 ( .A(B[8]), .B(\carry[0] ), .Y(\B_AS[8] ) );
  xor2a1 U3 ( .A(B[7]), .B(\carry[0] ), .Y(\B_AS[7] ) );
  xor2a1 U4 ( .A(B[6]), .B(\carry[0] ), .Y(\B_AS[6] ) );
  xor2a1 U5 ( .A(B[5]), .B(\carry[0] ), .Y(\B_AS[5] ) );
  xor2a1 U6 ( .A(B[4]), .B(\carry[0] ), .Y(\B_AS[4] ) );
  xor2a1 U7 ( .A(B[3]), .B(\carry[0] ), .Y(\B_AS[3] ) );
  xor2a1 U8 ( .A(B[2]), .B(\carry[0] ), .Y(\B_AS[2] ) );
  xor2a1 U9 ( .A(B[28]), .B(\carry[0] ), .Y(\B_AS[28] ) );
  xor2a1 U10 ( .A(B[27]), .B(\carry[0] ), .Y(\B_AS[27] ) );
  xor2a1 U11 ( .A(B[26]), .B(\carry[0] ), .Y(\B_AS[26] ) );
  xor2a1 U12 ( .A(B[25]), .B(\carry[0] ), .Y(\B_AS[25] ) );
  xor2a1 U13 ( .A(B[24]), .B(\carry[0] ), .Y(\B_AS[24] ) );
  xor2a1 U14 ( .A(B[23]), .B(\carry[0] ), .Y(\B_AS[23] ) );
  xor2a1 U15 ( .A(B[22]), .B(\carry[0] ), .Y(\B_AS[22] ) );
  xor2a1 U16 ( .A(B[21]), .B(\carry[0] ), .Y(\B_AS[21] ) );
  xor2a1 U17 ( .A(B[20]), .B(\carry[0] ), .Y(\B_AS[20] ) );
  xor2a1 U18 ( .A(B[1]), .B(\carry[0] ), .Y(\B_AS[1] ) );
  xor2a1 U19 ( .A(B[19]), .B(\carry[0] ), .Y(\B_AS[19] ) );
  xor2a1 U20 ( .A(B[18]), .B(\carry[0] ), .Y(\B_AS[18] ) );
  xor2a1 U21 ( .A(B[17]), .B(\carry[0] ), .Y(\B_AS[17] ) );
  xor2a1 U22 ( .A(B[16]), .B(\carry[0] ), .Y(\B_AS[16] ) );
  xor2a1 U23 ( .A(B[15]), .B(\carry[0] ), .Y(\B_AS[15] ) );
  xor2a1 U24 ( .A(B[14]), .B(\carry[0] ), .Y(\B_AS[14] ) );
  xor2a1 U25 ( .A(B[13]), .B(\carry[0] ), .Y(\B_AS[13] ) );
  xor2a1 U26 ( .A(B[12]), .B(\carry[0] ), .Y(\B_AS[12] ) );
  xor2a1 U27 ( .A(B[11]), .B(\carry[0] ), .Y(\B_AS[11] ) );
  xor2a1 U28 ( .A(B[10]), .B(\carry[0] ), .Y(\B_AS[10] ) );
  xor2a1 U29 ( .A(B[0]), .B(\carry[0] ), .Y(\B_AS[0] ) );
endmodule


module b14_DW01_addsub_0 ( A, B, CI, ADD_SUB, SUM, CO );
  input [28:0] A;
  input [28:0] B;
  output [28:0] SUM;
  input CI, ADD_SUB;
  output CO;
  wire   \carry[28] , \carry[27] , \carry[26] , \carry[25] , \carry[24] ,
         \carry[23] , \carry[22] , \carry[21] , \carry[20] , \carry[19] ,
         \carry[18] , \carry[17] , \carry[16] , \carry[15] , \carry[14] ,
         \carry[13] , \carry[12] , \carry[11] , \carry[10] , \carry[9] ,
         \carry[8] , \carry[7] , \carry[6] , \carry[5] , \carry[4] ,
         \carry[3] , \carry[2] , \carry[1] , \carry[0] , \B_AS[28] ,
         \B_AS[27] , \B_AS[26] , \B_AS[25] , \B_AS[24] , \B_AS[23] ,
         \B_AS[22] , \B_AS[21] , \B_AS[20] , \B_AS[19] , \B_AS[18] ,
         \B_AS[17] , \B_AS[16] , \B_AS[15] , \B_AS[14] , \B_AS[13] ,
         \B_AS[12] , \B_AS[11] , \B_AS[10] , \B_AS[9] , \B_AS[8] , \B_AS[7] ,
         \B_AS[6] , \B_AS[5] , \B_AS[4] , \B_AS[3] , \B_AS[2] , \B_AS[1] ,
         \B_AS[0] ;
  assign \carry[0]  = ADD_SUB;

  xor3a1 U1_28 ( .A(A[28]), .B(\B_AS[28] ), .C(\carry[28] ), .Y(SUM[28]) );
  fa1a1 U1_22 ( .A(A[22]), .B(\B_AS[22] ), .CI(\carry[22] ), .CO(\carry[23] ), 
        .S(SUM[22]) );
  fa1a1 U1_23 ( .A(A[23]), .B(\B_AS[23] ), .CI(\carry[23] ), .CO(\carry[24] ), 
        .S(SUM[23]) );
  fa1a1 U1_26 ( .A(A[26]), .B(\B_AS[26] ), .CI(\carry[26] ), .CO(\carry[27] ), 
        .S(SUM[26]) );
  fa1a1 U1_27 ( .A(A[27]), .B(\B_AS[27] ), .CI(\carry[27] ), .CO(\carry[28] ), 
        .S(SUM[27]) );
  fa1a1 U1_19 ( .A(A[19]), .B(\B_AS[19] ), .CI(\carry[19] ), .CO(\carry[20] ), 
        .S(SUM[19]) );
  fa1a1 U1_20 ( .A(A[20]), .B(\B_AS[20] ), .CI(\carry[20] ), .CO(\carry[21] ), 
        .S(SUM[20]) );
  fa1a1 U1_21 ( .A(A[21]), .B(\B_AS[21] ), .CI(\carry[21] ), .CO(\carry[22] ), 
        .S(SUM[21]) );
  fa1a1 U1_24 ( .A(A[24]), .B(\B_AS[24] ), .CI(\carry[24] ), .CO(\carry[25] ), 
        .S(SUM[24]) );
  fa1a1 U1_25 ( .A(A[25]), .B(\B_AS[25] ), .CI(\carry[25] ), .CO(\carry[26] ), 
        .S(SUM[25]) );
  fa1a1 U1_2 ( .A(A[2]), .B(\B_AS[2] ), .CI(\carry[2] ), .CO(\carry[3] ), .S(
        SUM[2]) );
  fa1a1 U1_3 ( .A(A[3]), .B(\B_AS[3] ), .CI(\carry[3] ), .CO(\carry[4] ), .S(
        SUM[3]) );
  fa1a1 U1_6 ( .A(A[6]), .B(\B_AS[6] ), .CI(\carry[6] ), .CO(\carry[7] ), .S(
        SUM[6]) );
  fa1a1 U1_7 ( .A(A[7]), .B(\B_AS[7] ), .CI(\carry[7] ), .CO(\carry[8] ), .S(
        SUM[7]) );
  fa1a1 U1_10 ( .A(A[10]), .B(\B_AS[10] ), .CI(\carry[10] ), .CO(\carry[11] ), 
        .S(SUM[10]) );
  fa1a1 U1_11 ( .A(A[11]), .B(\B_AS[11] ), .CI(\carry[11] ), .CO(\carry[12] ), 
        .S(SUM[11]) );
  fa1a1 U1_14 ( .A(A[14]), .B(\B_AS[14] ), .CI(\carry[14] ), .CO(\carry[15] ), 
        .S(SUM[14]) );
  fa1a1 U1_15 ( .A(A[15]), .B(\B_AS[15] ), .CI(\carry[15] ), .CO(\carry[16] ), 
        .S(SUM[15]) );
  fa1a1 U1_18 ( .A(A[18]), .B(\B_AS[18] ), .CI(\carry[18] ), .CO(\carry[19] ), 
        .S(SUM[18]) );
  fa1a1 U1_4 ( .A(A[4]), .B(\B_AS[4] ), .CI(\carry[4] ), .CO(\carry[5] ), .S(
        SUM[4]) );
  fa1a1 U1_5 ( .A(A[5]), .B(\B_AS[5] ), .CI(\carry[5] ), .CO(\carry[6] ), .S(
        SUM[5]) );
  fa1a1 U1_8 ( .A(A[8]), .B(\B_AS[8] ), .CI(\carry[8] ), .CO(\carry[9] ), .S(
        SUM[8]) );
  fa1a1 U1_9 ( .A(A[9]), .B(\B_AS[9] ), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  fa1a1 U1_12 ( .A(A[12]), .B(\B_AS[12] ), .CI(\carry[12] ), .CO(\carry[13] ), 
        .S(SUM[12]) );
  fa1a1 U1_13 ( .A(A[13]), .B(\B_AS[13] ), .CI(\carry[13] ), .CO(\carry[14] ), 
        .S(SUM[13]) );
  fa1a1 U1_16 ( .A(A[16]), .B(\B_AS[16] ), .CI(\carry[16] ), .CO(\carry[17] ), 
        .S(SUM[16]) );
  fa1a1 U1_17 ( .A(A[17]), .B(\B_AS[17] ), .CI(\carry[17] ), .CO(\carry[18] ), 
        .S(SUM[17]) );
  fa1a1 U1_1 ( .A(A[1]), .B(\B_AS[1] ), .CI(\carry[1] ), .CO(\carry[2] ), .S(
        SUM[1]) );
  fa1a1 U1_0 ( .A(A[0]), .B(\B_AS[0] ), .CI(\carry[0] ), .CO(\carry[1] ), .S(
        SUM[0]) );
  xor2a1 U1 ( .A(B[9]), .B(\carry[0] ), .Y(\B_AS[9] ) );
  xor2a1 U2 ( .A(B[8]), .B(\carry[0] ), .Y(\B_AS[8] ) );
  xor2a1 U3 ( .A(B[7]), .B(\carry[0] ), .Y(\B_AS[7] ) );
  xor2a1 U4 ( .A(B[6]), .B(\carry[0] ), .Y(\B_AS[6] ) );
  xor2a1 U5 ( .A(B[5]), .B(\carry[0] ), .Y(\B_AS[5] ) );
  xor2a1 U6 ( .A(B[4]), .B(\carry[0] ), .Y(\B_AS[4] ) );
  xor2a1 U7 ( .A(B[3]), .B(\carry[0] ), .Y(\B_AS[3] ) );
  xor2a1 U8 ( .A(B[2]), .B(\carry[0] ), .Y(\B_AS[2] ) );
  xor2a1 U9 ( .A(B[28]), .B(\carry[0] ), .Y(\B_AS[28] ) );
  xor2a1 U10 ( .A(B[27]), .B(\carry[0] ), .Y(\B_AS[27] ) );
  xor2a1 U11 ( .A(B[26]), .B(\carry[0] ), .Y(\B_AS[26] ) );
  xor2a1 U12 ( .A(B[25]), .B(\carry[0] ), .Y(\B_AS[25] ) );
  xor2a1 U13 ( .A(B[24]), .B(\carry[0] ), .Y(\B_AS[24] ) );
  xor2a1 U14 ( .A(B[23]), .B(\carry[0] ), .Y(\B_AS[23] ) );
  xor2a1 U15 ( .A(B[22]), .B(\carry[0] ), .Y(\B_AS[22] ) );
  xor2a1 U16 ( .A(B[21]), .B(\carry[0] ), .Y(\B_AS[21] ) );
  xor2a1 U17 ( .A(B[20]), .B(\carry[0] ), .Y(\B_AS[20] ) );
  xor2a1 U18 ( .A(B[1]), .B(\carry[0] ), .Y(\B_AS[1] ) );
  xor2a1 U19 ( .A(B[19]), .B(\carry[0] ), .Y(\B_AS[19] ) );
  xor2a1 U20 ( .A(B[18]), .B(\carry[0] ), .Y(\B_AS[18] ) );
  xor2a1 U21 ( .A(B[17]), .B(\carry[0] ), .Y(\B_AS[17] ) );
  xor2a1 U22 ( .A(B[16]), .B(\carry[0] ), .Y(\B_AS[16] ) );
  xor2a1 U23 ( .A(B[15]), .B(\carry[0] ), .Y(\B_AS[15] ) );
  xor2a1 U24 ( .A(B[14]), .B(\carry[0] ), .Y(\B_AS[14] ) );
  xor2a1 U25 ( .A(B[13]), .B(\carry[0] ), .Y(\B_AS[13] ) );
  xor2a1 U26 ( .A(B[12]), .B(\carry[0] ), .Y(\B_AS[12] ) );
  xor2a1 U27 ( .A(B[11]), .B(\carry[0] ), .Y(\B_AS[11] ) );
  xor2a1 U28 ( .A(B[10]), .B(\carry[0] ), .Y(\B_AS[10] ) );
  xor2a1 U29 ( .A(B[0]), .B(\carry[0] ), .Y(\B_AS[0] ) );
endmodule


module b14 ( clock, reset, .addr({\addr[19] , \addr[18] , \addr[17] , 
        \addr[16] , \addr[15] , \addr[14] , \addr[13] , \addr[12] , \addr[11] , 
        \addr[10] , \addr[9] , \addr[8] , \addr[7] , \addr[6] , \addr[5] , 
        \addr[4] , \addr[3] , \addr[2] , \addr[1] , \addr[0] }), .datai({
        \datai[31] , \datai[30] , \datai[29] , \datai[28] , \datai[27] , 
        \datai[26] , \datai[25] , \datai[24] , \datai[23] , \datai[22] , 
        \datai[21] , \datai[20] , \datai[19] , \datai[18] , \datai[17] , 
        \datai[16] , \datai[15] , \datai[14] , \datai[13] , \datai[12] , 
        \datai[11] , \datai[10] , \datai[9] , \datai[8] , \datai[7] , 
        \datai[6] , \datai[5] , \datai[4] , \datai[3] , \datai[2] , \datai[1] , 
        \datai[0] }), .datao({\datao[31] , \datao[30] , \datao[29] , 
        \datao[28] , \datao[27] , \datao[26] , \datao[25] , \datao[24] , 
        \datao[23] , \datao[22] , \datao[21] , \datao[20] , \datao[19] , 
        \datao[18] , \datao[17] , \datao[16] , \datao[15] , \datao[14] , 
        \datao[13] , \datao[12] , \datao[11] , \datao[10] , \datao[9] , 
        \datao[8] , \datao[7] , \datao[6] , \datao[5] , \datao[4] , \datao[3] , 
        \datao[2] , \datao[1] , \datao[0] }), rd, wr );
  input clock, reset, \datai[31] , \datai[30] , \datai[29] , \datai[28] ,
         \datai[27] , \datai[26] , \datai[25] , \datai[24] , \datai[23] ,
         \datai[22] , \datai[21] , \datai[20] , \datai[19] , \datai[18] ,
         \datai[17] , \datai[16] , \datai[15] , \datai[14] , \datai[13] ,
         \datai[12] , \datai[11] , \datai[10] , \datai[9] , \datai[8] ,
         \datai[7] , \datai[6] , \datai[5] , \datai[4] , \datai[3] ,
         \datai[2] , \datai[1] , \datai[0] ;
  output \addr[19] , \addr[18] , \addr[17] , \addr[16] , \addr[15] ,
         \addr[14] , \addr[13] , \addr[12] , \addr[11] , \addr[10] , \addr[9] ,
         \addr[8] , \addr[7] , \addr[6] , \addr[5] , \addr[4] , \addr[3] ,
         \addr[2] , \addr[1] , \addr[0] , \datao[31] , \datao[30] ,
         \datao[29] , \datao[28] , \datao[27] , \datao[26] , \datao[25] ,
         \datao[24] , \datao[23] , \datao[22] , \datao[21] , \datao[20] ,
         \datao[19] , \datao[18] , \datao[17] , \datao[16] , \datao[15] ,
         \datao[14] , \datao[13] , \datao[12] , \datao[11] , \datao[10] ,
         \datao[9] , \datao[8] , \datao[7] , \datao[6] , \datao[5] ,
         \datao[4] , \datao[3] , \datao[2] , \datao[1] , \datao[0] , rd, wr;
  wire   B, state, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302,
         N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545,
         N546, N547, N548, N549, N550, N551, N552, N553, N554, N555, N556,
         N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567,
         N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578,
         N579, N580, N581, N582, N583, N584, N585, N654, N655, N656, N657,
         N658, N659, N660, N661, N662, N663, N664, N665, N666, N667, N668,
         N669, N670, N671, N672, N673, N674, N675, N676, N677, N678, N679,
         N680, N681, N682, N683, N684, N685, N847, N849, N939, N940, N941,
         N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952,
         N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963,
         N964, N965, N966, N967, N968, N969, N970, N1028, N1029, N1030, N1031,
         N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041,
         N1042, N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051,
         N1052, N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1315, N1316,
         N1317, N1318, N1319, N1320, N1321, N1322, N1323, N1324, N1325, N1326,
         N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1336,
         N1337, N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346,
         N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354, N2117, N2118,
         N2119, N2120, N2121, N2122, N2123, N2124, N2125, N2126, N2127, N2128,
         N2129, N2130, N2131, N2132, N2133, N2134, N2135, N2136, N2137, N2138,
         N2139, N2140, N2141, N2142, N2143, N2144, N2145, N2146, N2525, N2526,
         N2527, N2528, N2529, N2530, N2531, N2532, N2533, N2534, N2535, N2536,
         N2537, N2538, N2539, N2540, N2541, N2542, N2543, N2544, N2545, N2546,
         N2547, N2548, N2549, N2550, N2551, N2552, N2553, N2554, N2933, N2934,
         N2935, N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2943, N2944,
         N2945, N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954,
         N2955, N2956, N2957, N2958, N2959, N2960, N2961, N2962, N3341, N3342,
         N3343, N3344, N3345, N3346, N3347, N3348, N3349, N3350, N3351, N3352,
         N3353, N3354, N3355, N3356, N3357, N3358, N3359, N3360, N3361, N3362,
         N3363, N3364, N3365, N3366, N3367, N3368, N3369, N3370, N3749, N3750,
         N3751, N3752, N3753, N3754, N3755, N3756, N3757, N3758, N3759, N3760,
         N3761, N3762, N3763, N3764, N3765, N3766, N3767, N3768, N3769, N3770,
         N3771, N3772, N3773, N3774, N3775, N3776, N3777, N3778, N4157, N4158,
         N4159, N4160, N4161, N4162, N4163, N4164, N4165, N4166, N4167, N4168,
         N4169, N4170, N4171, N4172, N4173, N4174, N4175, N4176, N4177, N4178,
         N4179, N4180, N4181, N4182, N4183, N4184, N4185, N4186, N4565, N4566,
         N4567, N4568, N4569, N4570, N4571, N4572, N4573, N4574, N4575, N4576,
         N4577, N4578, N4579, N4580, N4581, N4582, N4583, N4584, N4585, N4586,
         N4587, N4588, N4589, N4590, N4591, N4592, N4593, N4594, N4655, N4656,
         N4657, N4658, N4659, N4660, N4661, N4662, N4663, N4664, N4665, N4666,
         N4667, N4668, N4669, N4670, N4671, N4672, N4673, N4674, N4675, N4676,
         N4677, N4678, N4679, N4680, N4681, N4682, N4683, N4973, N4974, N4975,
         N4976, N4977, N4978, N4979, N4980, N4981, N4982, N4983, N4984, N4985,
         N4986, N4987, N4988, N4989, N4990, N4991, N4992, N4993, N4994, N4995,
         N4996, N4997, N4998, N4999, N5000, N5001, N5002, N5654, N5656, N5658,
         N5660, N5662, N5664, N5666, N5668, N5670, N5672, N5674, N5676, N5678,
         N5680, N5682, N5684, N5686, N5688, N5690, N5692, N5694, N5696, N5698,
         N5700, N5702, N5704, N5706, N5708, N5710, N5712, N5718, N5720, N5722,
         N5724, N5726, N5728, N5730, N5732, N5734, N5736, N5738, N5740, N5742,
         N5744, N5746, N5748, N5750, N5752, N5754, N5756, N5758, N5760, N5762,
         N5764, N5766, N5768, N5770, N5772, N5774, N5776, N5778, N5780, N6175,
         N6305, N6717, N6754, N6892, N6893, N6894, N6895, N6896, N6897, N6898,
         N6899, N6900, N6901, N6902, N6903, N6904, N6905, N6906, N6907, N6908,
         N6909, N6910, N6911, N6912, N6913, N6914, N6915, N6916, N6917, N6918,
         N6919, N6920, N6954, N6956, N6958, N6960, N6962, N6964, N6966, N6968,
         N6970, N6972, N6974, N6976, N6978, N6980, N6982, N6984, N6986, N6988,
         N6990, N6991, N6992, N6993, N6995, N6997, N6999, N7001, N7003, N7005,
         N7007, N7009, N7011, N7013, N7015, N7017, N7019, N7021, N7023, N7025,
         N7027, N7029, N7031, N7033, N7035, N7037, N7039, N7041, N7043, N7045,
         N7047, N7049, N7051, N7053, N7055, N7056, N7057, N7058, N7091, N7123,
         N7124, N7156, N7188, N7220, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, \U3/U1/Z_0 , \U3/U1/Z_1 , \U3/U1/Z_2 ,
         \U3/U1/Z_3 , \U3/U1/Z_4 , \U3/U1/Z_5 , \U3/U1/Z_6 , \U3/U1/Z_7 ,
         \U3/U1/Z_8 , \U3/U1/Z_9 , \U3/U1/Z_10 , \U3/U1/Z_11 , \U3/U1/Z_12 ,
         \U3/U1/Z_13 , \U3/U1/Z_14 , \U3/U1/Z_15 , \U3/U1/Z_16 , \U3/U1/Z_17 ,
         \U3/U1/Z_18 , \U3/U1/Z_19 , \U3/U1/Z_20 , \U3/U1/Z_21 , \U3/U1/Z_22 ,
         \U3/U1/Z_23 , \U3/U1/Z_24 , \U3/U1/Z_25 , \U3/U1/Z_26 , \U3/U1/Z_27 ,
         \U3/U1/Z_28 , \U3/U2/Z_0 , \U3/U3/Z_0 , \U3/U3/Z_1 , \U3/U3/Z_2 ,
         \U3/U3/Z_3 , \U3/U3/Z_4 , \U3/U3/Z_5 , \U3/U3/Z_6 , \U3/U3/Z_7 ,
         \U3/U3/Z_8 , \U3/U3/Z_9 , \U3/U3/Z_10 , \U3/U3/Z_11 , \U3/U3/Z_12 ,
         \U3/U3/Z_13 , \U3/U3/Z_14 , \U3/U3/Z_15 , \U3/U3/Z_16 , \U3/U3/Z_17 ,
         \U3/U3/Z_18 , \U3/U3/Z_19 , \U3/U3/Z_20 , \U3/U3/Z_21 , \U3/U3/Z_22 ,
         \U3/U3/Z_23 , \U3/U3/Z_24 , \U3/U3/Z_25 , \U3/U3/Z_26 , \U3/U3/Z_27 ,
         \U3/U3/Z_28 , \U3/U4/Z_0 , \U3/U4/Z_1 , \U3/U4/Z_2 , \U3/U4/Z_3 ,
         \U3/U4/Z_4 , \U3/U4/Z_5 , \U3/U4/Z_6 , \U3/U4/Z_7 , \U3/U4/Z_8 ,
         \U3/U4/Z_9 , \U3/U4/Z_10 , \U3/U4/Z_11 , \U3/U4/Z_12 , \U3/U4/Z_13 ,
         \U3/U4/Z_14 , \U3/U4/Z_15 , \U3/U4/Z_16 , \U3/U4/Z_17 , \U3/U4/Z_18 ,
         \U3/U4/Z_19 , \U3/U4/Z_20 , \U3/U4/Z_21 , \U3/U4/Z_22 , \U3/U4/Z_23 ,
         \U3/U4/Z_24 , \U3/U4/Z_25 , \U3/U4/Z_26 , \U3/U4/Z_27 , \U3/U4/Z_28 ,
         \U3/U5/Z_0 , \U3/U6/Z_0 , \U3/U6/Z_1 , \U3/U6/Z_2 , \U3/U6/Z_3 ,
         \U3/U6/Z_4 , \U3/U6/Z_5 , \U3/U6/Z_6 , \U3/U6/Z_7 , \U3/U6/Z_8 ,
         \U3/U6/Z_9 , \U3/U6/Z_10 , \U3/U6/Z_11 , \U3/U6/Z_12 , \U3/U6/Z_13 ,
         \U3/U6/Z_14 , \U3/U6/Z_15 , \U3/U6/Z_16 , \U3/U6/Z_17 , \U3/U6/Z_18 ,
         \U3/U6/Z_19 , \U3/U6/Z_20 , \U3/U6/Z_21 , \U3/U6/Z_22 , \U3/U6/Z_23 ,
         \U3/U6/Z_24 , \U3/U6/Z_25 , \U3/U6/Z_26 , \U3/U6/Z_27 , \U3/U6/Z_28 ,
         \U3/U6/Z_29 , \U3/U6/Z_30 , \U3/U6/Z_31 , \U3/U7/Z_0 , \U3/U7/Z_1 ,
         \U3/U7/Z_2 , \U3/U7/Z_3 , \U3/U7/Z_4 , \U3/U7/Z_5 , \U3/U7/Z_6 ,
         \U3/U7/Z_7 , \U3/U7/Z_8 , \U3/U7/Z_9 , \U3/U7/Z_10 , \U3/U7/Z_11 ,
         \U3/U7/Z_12 , \U3/U7/Z_13 , \U3/U7/Z_14 , \U3/U7/Z_15 , \U3/U7/Z_16 ,
         \U3/U7/Z_17 , \U3/U7/Z_18 , \U3/U7/Z_19 , \U3/U7/Z_20 , \U3/U7/Z_21 ,
         \U3/U7/Z_22 , \U3/U7/Z_23 , \U3/U7/Z_24 , \U3/U7/Z_25 , \U3/U7/Z_26 ,
         \U3/U7/Z_27 , \U3/U7/Z_28 , \U3/U7/Z_29 , \U3/U7/Z_30 , \U3/U7/Z_31 ,
         \U3/U8/Z_0 , \U3/U8/Z_1 , \U3/U8/Z_2 , \U3/U8/Z_3 , \U3/U8/Z_4 ,
         \U3/U8/Z_5 , \U3/U8/Z_6 , \U3/U8/Z_7 , \U3/U8/Z_8 , \U3/U8/Z_9 ,
         \U3/U8/Z_10 , \U3/U8/Z_11 , \U3/U8/Z_12 , \U3/U8/Z_13 , \U3/U8/Z_14 ,
         \U3/U8/Z_15 , \U3/U8/Z_16 , \U3/U8/Z_17 , \U3/U8/Z_18 , \U3/U8/Z_19 ,
         \U3/U8/Z_20 , \U3/U8/Z_21 , \U3/U8/Z_22 , \U3/U8/Z_23 , \U3/U8/Z_24 ,
         \U3/U8/Z_25 , \U3/U8/Z_26 , \U3/U8/Z_27 , \U3/U8/Z_28 , \U3/U8/Z_29 ,
         \U3/U8/Z_30 , \U3/U8/Z_31 , \U3/U9/Z_0 , \U3/U9/Z_1 , \U3/U9/Z_2 ,
         \U3/U9/Z_3 , \U3/U9/Z_4 , \U3/U9/Z_5 , \U3/U9/Z_6 , \U3/U9/Z_7 ,
         \U3/U9/Z_8 , \U3/U9/Z_9 , \U3/U9/Z_10 , \U3/U9/Z_11 , \U3/U9/Z_12 ,
         \U3/U9/Z_13 , \U3/U9/Z_14 , \U3/U9/Z_15 , \U3/U9/Z_16 , \U3/U9/Z_17 ,
         \U3/U9/Z_18 , \U3/U9/Z_30 , \U3/U9/Z_31 , \U3/U10/Z_0 , n425, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745;
  wire   [31:0] IR;
  wire   [31:0] d;
  wire   [31:0] reg0;
  wire   [31:0] reg1;
  wire   [31:0] reg2;
  wire   [28:0] reg3;
  wire   SYNOPSYS_UNCONNECTED__0;

  b14_DW01_addsub_0 r798 ( .A({N682, N681, N680, N679, N678, N677, N676, N675, 
        N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, 
        N662, N661, N660, N659, N658, N657, N656, N655, N654}), .B({
        \U3/U1/Z_28 , \U3/U1/Z_27 , \U3/U1/Z_26 , \U3/U1/Z_25 , \U3/U1/Z_24 , 
        \U3/U1/Z_23 , \U3/U1/Z_22 , \U3/U1/Z_21 , \U3/U1/Z_20 , \U3/U1/Z_19 , 
        \U3/U1/Z_18 , \U3/U1/Z_17 , \U3/U1/Z_16 , \U3/U1/Z_15 , \U3/U1/Z_14 , 
        \U3/U1/Z_13 , \U3/U1/Z_12 , \U3/U1/Z_11 , \U3/U1/Z_10 , \U3/U1/Z_9 , 
        \U3/U1/Z_8 , \U3/U1/Z_7 , \U3/U1/Z_6 , \U3/U1/Z_5 , \U3/U1/Z_4 , 
        \U3/U1/Z_3 , \U3/U1/Z_2 , \U3/U1/Z_1 , \U3/U1/Z_0 }), .CI(0), 
        .ADD_SUB(\U3/U2/Z_0 ), .SUM({N4683, N4682, N4681, N4680, N4679, N4678, 
        N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, 
        N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659, N4658, 
        N4657, N4656, N4655}) );
  b14_DW01_addsub_1 r794 ( .A({\U3/U3/Z_28 , \U3/U3/Z_27 , \U3/U3/Z_26 , 
        \U3/U3/Z_25 , \U3/U3/Z_24 , \U3/U3/Z_23 , \U3/U3/Z_22 , \U3/U3/Z_21 , 
        \U3/U3/Z_20 , \U3/U3/Z_19 , \U3/U3/Z_18 , \U3/U3/Z_17 , \U3/U3/Z_16 , 
        \U3/U3/Z_15 , \U3/U3/Z_14 , \U3/U3/Z_13 , \U3/U3/Z_12 , \U3/U3/Z_11 , 
        \U3/U3/Z_10 , \U3/U3/Z_9 , \U3/U3/Z_8 , \U3/U3/Z_7 , \U3/U3/Z_6 , 
        \U3/U3/Z_5 , \U3/U3/Z_4 , \U3/U3/Z_3 , \U3/U3/Z_2 , \U3/U3/Z_1 , 
        \U3/U3/Z_0 }), .B({\U3/U4/Z_28 , \U3/U4/Z_27 , \U3/U4/Z_26 , 
        \U3/U4/Z_25 , \U3/U4/Z_24 , \U3/U4/Z_23 , \U3/U4/Z_22 , \U3/U4/Z_21 , 
        \U3/U4/Z_20 , \U3/U4/Z_19 , \U3/U4/Z_18 , \U3/U4/Z_17 , \U3/U4/Z_16 , 
        \U3/U4/Z_15 , \U3/U4/Z_14 , \U3/U4/Z_13 , \U3/U4/Z_12 , \U3/U4/Z_11 , 
        \U3/U4/Z_10 , \U3/U4/Z_9 , \U3/U4/Z_8 , \U3/U4/Z_7 , \U3/U4/Z_6 , 
        \U3/U4/Z_5 , \U3/U4/Z_4 , \U3/U4/Z_3 , \U3/U4/Z_2 , \U3/U4/Z_1 , 
        \U3/U4/Z_0 }), .CI(0), .ADD_SUB(\U3/U5/Z_0 ), .SUM({n33, n34, n35, 
        n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
        n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61}) );
  b14_DW01_cmp2_0 r795 ( .A({\U3/U6/Z_31 , \U3/U6/Z_30 , \U3/U6/Z_29 , 
        \U3/U6/Z_28 , \U3/U6/Z_27 , \U3/U6/Z_26 , \U3/U6/Z_25 , \U3/U6/Z_24 , 
        \U3/U6/Z_23 , \U3/U6/Z_22 , \U3/U6/Z_21 , \U3/U6/Z_20 , \U3/U6/Z_19 , 
        \U3/U6/Z_18 , \U3/U6/Z_17 , \U3/U6/Z_16 , \U3/U6/Z_15 , \U3/U6/Z_14 , 
        \U3/U6/Z_13 , \U3/U6/Z_12 , \U3/U6/Z_11 , \U3/U6/Z_10 , \U3/U6/Z_9 , 
        \U3/U6/Z_8 , \U3/U6/Z_7 , \U3/U6/Z_6 , \U3/U6/Z_5 , \U3/U6/Z_4 , 
        \U3/U6/Z_3 , \U3/U6/Z_2 , \U3/U6/Z_1 , \U3/U6/Z_0 }), .B({\U3/U7/Z_31 , 
        \U3/U7/Z_30 , \U3/U7/Z_29 , \U3/U7/Z_28 , \U3/U7/Z_27 , \U3/U7/Z_26 , 
        \U3/U7/Z_25 , \U3/U7/Z_24 , \U3/U7/Z_23 , \U3/U7/Z_22 , \U3/U7/Z_21 , 
        \U3/U7/Z_20 , \U3/U7/Z_19 , \U3/U7/Z_18 , \U3/U7/Z_17 , \U3/U7/Z_16 , 
        \U3/U7/Z_15 , \U3/U7/Z_14 , \U3/U7/Z_13 , \U3/U7/Z_12 , \U3/U7/Z_11 , 
        \U3/U7/Z_10 , \U3/U7/Z_9 , \U3/U7/Z_8 , \U3/U7/Z_7 , \U3/U7/Z_6 , 
        \U3/U7/Z_5 , \U3/U7/Z_4 , \U3/U7/Z_3 , \U3/U7/Z_2 , \U3/U7/Z_1 , 
        \U3/U7/Z_0 }), .LEQ(0), .TC(1), .LT_LE(N6717) );
  b14_DW01_addsub_2 r796 ( .A({\U3/U8/Z_31 , \U3/U8/Z_30 , \U3/U8/Z_29 , 
        \U3/U8/Z_28 , \U3/U8/Z_27 , \U3/U8/Z_26 , \U3/U8/Z_25 , \U3/U8/Z_24 , 
        \U3/U8/Z_23 , \U3/U8/Z_22 , \U3/U8/Z_21 , \U3/U8/Z_20 , \U3/U8/Z_19 , 
        \U3/U8/Z_18 , \U3/U8/Z_17 , \U3/U8/Z_16 , \U3/U8/Z_15 , \U3/U8/Z_14 , 
        \U3/U8/Z_13 , \U3/U8/Z_12 , \U3/U8/Z_11 , \U3/U8/Z_10 , \U3/U8/Z_9 , 
        \U3/U8/Z_8 , \U3/U8/Z_7 , \U3/U8/Z_6 , \U3/U8/Z_5 , \U3/U8/Z_4 , 
        \U3/U8/Z_3 , \U3/U8/Z_2 , \U3/U8/Z_1 , \U3/U8/Z_0 }), .B({\U3/U9/Z_31 , 
        \U3/U9/Z_30 , \U3/U9/Z_31 , \U3/U9/Z_31 , \U3/U9/Z_31 , \U3/U9/Z_31 , 
        \U3/U9/Z_31 , \U3/U9/Z_31 , \U3/U9/Z_31 , \U3/U9/Z_31 , \U3/U9/Z_31 , 
        \U3/U9/Z_31 , \U3/U9/Z_31 , \U3/U9/Z_18 , \U3/U9/Z_17 , \U3/U9/Z_16 , 
        \U3/U9/Z_15 , \U3/U9/Z_14 , \U3/U9/Z_13 , \U3/U9/Z_12 , \U3/U9/Z_11 , 
        \U3/U9/Z_10 , \U3/U9/Z_9 , \U3/U9/Z_8 , \U3/U9/Z_7 , \U3/U9/Z_6 , 
        \U3/U9/Z_5 , \U3/U9/Z_4 , \U3/U9/Z_3 , \U3/U9/Z_2 , \U3/U9/Z_1 , 
        \U3/U9/Z_0 }), .CI(0), .ADD_SUB(\U3/U10/Z_0 ), .SUM({n189, n190, 
        n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
        n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
        n215, n216, n217, n218, n219, n220}) );
  b14_DW01_cmp6_0 r620 ( .A({N685, N684, N683, N682, N681, N680, N679, N678, 
        N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, 
        N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654}), .B({N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, 
        N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, 
        N946, N945, N944, N943, N942, N941, N940, N939}), .TC(1), .LT(N6175), .GT(N6305) );
  b14_DW01_sub_0 r612 ( .A({N683, N682, N681, N680, N679, N678, N677, N676, 
        N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, 
        N663, N662, N661, N660, N659, N658, N657, N656, N655, N654}), .B({N968, 
        N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, 
        N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, 
        N943, N942, N941, N940, N939}), .CI(0), .DIFF({N5002, N5001, N5000, 
        N4999, N4998, N4997, N4996, N4995, N4994, N4993, N4992, N4991, N4990, 
        N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, 
        N4979, N4978, N4977, N4976, N4975, N4974, N4973}) );
  b14_DW01_add_0 r608 ( .A({N683, N682, N681, N680, N679, N678, N677, N676, 
        N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, 
        N663, N662, N661, N660, N659, N658, N657, N656, N655, N654}), .B({N968, 
        N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, 
        N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, 
        N943, N942, N941, N940, N939}), .CI(0), .SUM({N4594, N4593, N4592, 
        N4591, N4590, N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582, 
        N4581, N4580, N4579, N4578, N4577, N4576, N4575, N4574, N4573, N4572, 
        N4571, N4570, N4569, N4568, N4567, N4566, N4565}) );
  b14_DW01_sub_1 r604 ( .A({N683, N682, N681, N680, N679, N678, N677, N676, 
        N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, 
        N663, N662, N661, N660, N659, N658, N657, N656, N655, N654}), .B({N968, 
        N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, 
        N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, 
        N943, N942, N941, N940, N939}), .CI(0), .DIFF({N4186, N4185, N4184, 
        N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, 
        N4173, N4172, N4171, N4170, N4169, N4168, N4167, N4166, N4165, N4164, 
        N4163, N4162, N4161, N4160, N4159, N4158, N4157}) );
  b14_DW01_add_1 r600 ( .A({N683, N682, N681, N680, N679, N678, N677, N676, 
        N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, 
        N663, N662, N661, N660, N659, N658, N657, N656, N655, N654}), .B({N968, 
        N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, 
        N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, 
        N943, N942, N941, N940, N939}), .CI(0), .SUM({N3778, N3777, N3776, 
        N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, 
        N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, 
        N3755, N3754, N3753, N3752, N3751, N3750, N3749}) );
  b14_DW01_sub_2 r596 ( .A({N683, N682, N681, N680, N679, N678, N677, N676, 
        N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, 
        N663, N662, N661, N660, N659, N658, N657, N656, N655, N654}), .B({N968, 
        N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, 
        N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, 
        N943, N942, N941, N940, N939}), .CI(0), .DIFF({N3370, N3369, N3368, 
        N3367, N3366, N3365, N3364, N3363, N3362, N3361, N3360, N3359, N3358, 
        N3357, N3356, N3355, N3354, N3353, N3352, N3351, N3350, N3349, N3348, 
        N3347, N3346, N3345, N3344, N3343, N3342, N3341}) );
  b14_DW01_sub_3 r592 ( .A({N683, N682, N681, N680, N679, N678, N677, N676, 
        N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, 
        N663, N662, N661, N660, N659, N658, N657, N656, N655, N654}), .B({N968, 
        N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, 
        N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, 
        N943, N942, N941, N940, N939}), .CI(0), .DIFF({N2962, N2961, N2960, 
        N2959, N2958, N2957, N2956, N2955, N2954, N2953, N2952, N2951, N2950, 
        N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, 
        N2939, N2938, N2937, N2936, N2935, N2934, N2933}) );
  b14_DW01_add_2 r588 ( .A({N683, N682, N681, N680, N679, N678, N677, N676, 
        N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, 
        N663, N662, N661, N660, N659, N658, N657, N656, N655, N654}), .B({N968, 
        N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, 
        N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, 
        N943, N942, N941, N940, N939}), .CI(0), .SUM({N2554, N2553, N2552, 
        N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, 
        N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, 
        N2531, N2530, N2529, N2528, N2527, N2526, N2525}) );
  b14_DW01_add_3 r584 ( .A({N683, N682, N681, N680, N679, N678, N677, N676, 
        N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, 
        N663, N662, N661, N660, N659, N658, N657, N656, N655, N654}), .B({N968, 
        N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, 
        N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, 
        N943, N942, N941, N940, N939}), .CI(0), .SUM({N2146, N2145, N2144, 
        N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, 
        N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, 
        N2123, N2122, N2121, N2120, N2119, N2118, N2117}) );
  b14_DW01_add_4 r581 ( .A({N536, N537, N538, N539, N540, N541, N542, N543, 
        N544, N545, N546, N547, N548, N549, N550, N551, N552, N553, N554, N555}), .B(reg2[19:0]), .CI(0), .SUM({N1354, N1353, N1352, N1351, N1350, N1349, 
        N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, 
        N1338, N1337, N1336, N1335}) );
  b14_DW01_add_5 r580 ( .A({N536, N537, N538, N539, N540, N541, N542, N543, 
        N544, N545, N546, N547, N548, N549, N550, N551, N552, N553, N554, N555}), .B(reg1[19:0]), .CI(0), .SUM({N1334, N1333, N1332, N1331, N1330, N1329, 
        N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, 
        N1318, N1317, N1316, N1315}) );
  b14_DW01_sub_4 r578 ( .A({0, 0, 0, 0, 0, 0, 0, 0, 
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}), .B({N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, 
        N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, 
        N946, N945, N944, N943, N942, N941, N940, N939}), .CI(0), .DIFF({
        N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, 
        N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, 
        N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, 
        N1029, N1028}) );
  b14_DW01_sub_5 sub_84 ( .A({0, 0, 0, 0, 0, 0, 0, 0, 
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}), .B({N325, IR[30:0]}), .CI(0), .DIFF({N324, N323, N322, N321, N320, N319, 
        N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, 
        N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, 
        N294, N293}) );
  b14_DW01_add_7 add_95 ( .A({0, 0, reg3}), .B({0, 0, 0, 0, 
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
        0, 0, 0}), .CI(0), .SUM({SYNOPSYS_UNCONNECTED__0, N585, 
        N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, 
        N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, 
        N560, N559, N558, N557, N556}) );
  fdef2a6 \d_reg[1]  ( .D(N849), .E(N7123), .CLK(clock), .CLR(n2177), .Q(d[1])
         );
  fdef2a6 \d_reg[0]  ( .D(N847), .E(N7123), .CLK(clock), .CLR(n2177), .Q(d[0])
         );
  fdef2a6 \reg2_reg[20]  ( .D(N5758), .E(N7220), .CLK(clock), .CLR(n2156), .Q(
        reg2[20]) );
  fdef2a6 \reg2_reg[21]  ( .D(N5760), .E(N7220), .CLK(clock), .CLR(n2155), .Q(
        reg2[21]) );
  fdef2a6 \reg2_reg[22]  ( .D(N5762), .E(N7220), .CLK(clock), .CLR(n2154), .Q(
        reg2[22]) );
  fdef2a6 \reg2_reg[23]  ( .D(N5764), .E(N7220), .CLK(clock), .CLR(n2153), .Q(
        reg2[23]) );
  fdef2a6 \reg2_reg[24]  ( .D(N5766), .E(N7220), .CLK(clock), .CLR(n2152), .Q(
        reg2[24]) );
  fdef2a6 \reg2_reg[25]  ( .D(N5768), .E(N7220), .CLK(clock), .CLR(n2151), .Q(
        reg2[25]) );
  fdef2a6 \reg2_reg[26]  ( .D(N5770), .E(N7220), .CLK(clock), .CLR(n2150), .Q(
        reg2[26]) );
  fdef2a6 \reg2_reg[27]  ( .D(N5772), .E(N7220), .CLK(clock), .CLR(n2149), .Q(
        reg2[27]) );
  fdef2a6 \reg2_reg[28]  ( .D(N5774), .E(N7220), .CLK(clock), .CLR(n2148), .Q(
        reg2[28]) );
  fdef2a6 \reg2_reg[29]  ( .D(N5776), .E(N7220), .CLK(clock), .CLR(n2146), .Q(
        reg2[29]) );
  fdef2a6 \reg0_reg[29]  ( .D(N5712), .E(N7156), .CLK(clock), .CLR(n2146), .Q(
        reg0[29]) );
  fdef2a6 \reg0_reg[27]  ( .D(N5708), .E(N7156), .CLK(clock), .CLR(n2150), .Q(
        reg0[27]) );
  fdef2a6 \reg0_reg[25]  ( .D(N5704), .E(N7156), .CLK(clock), .CLR(n2152), .Q(
        reg0[25]) );
  fdef2a6 \reg0_reg[23]  ( .D(N5700), .E(N7156), .CLK(clock), .CLR(n2154), .Q(
        reg0[23]) );
  fdef2a6 \reg0_reg[21]  ( .D(N5696), .E(N7156), .CLK(clock), .CLR(n2156), .Q(
        reg0[21]) );
  fdef2a6 \reg0_reg[19]  ( .D(N5692), .E(N7156), .CLK(clock), .CLR(n2158), .Q(
        reg0[19]) );
  fdef2a6 \reg0_reg[17]  ( .D(N5688), .E(N7156), .CLK(clock), .CLR(n2160), .Q(
        reg0[17]) );
  fdef2a6 \reg0_reg[15]  ( .D(N5684), .E(N7156), .CLK(clock), .CLR(n2162), .Q(
        reg0[15]) );
  fdef2a6 \reg0_reg[13]  ( .D(N5680), .E(N7156), .CLK(clock), .CLR(n2164), .Q(
        reg0[13]) );
  fdef2a6 \reg0_reg[11]  ( .D(N5676), .E(N7156), .CLK(clock), .CLR(n2166), .Q(
        reg0[11]) );
  fdef2a6 \reg0_reg[9]  ( .D(N5672), .E(N7156), .CLK(clock), .CLR(n2168), .Q(
        reg0[9]) );
  fdef2a6 \reg0_reg[7]  ( .D(N5668), .E(N7156), .CLK(clock), .CLR(n2170), .Q(
        reg0[7]) );
  fdef2a6 \reg0_reg[5]  ( .D(N5664), .E(N7156), .CLK(clock), .CLR(n2172), .Q(
        reg0[5]) );
  fdef2a6 \reg0_reg[3]  ( .D(N5660), .E(N7156), .CLK(clock), .CLR(n2174), .Q(
        reg0[3]) );
  fdef2a6 \reg0_reg[1]  ( .D(N5656), .E(N7156), .CLK(clock), .CLR(n2176), .Q(
        reg0[1]) );
  fdef2a6 \reg0_reg[2]  ( .D(N5658), .E(N7156), .CLK(clock), .CLR(n2175), .Q(
        reg0[2]) );
  fdef2a6 \reg0_reg[4]  ( .D(N5662), .E(N7156), .CLK(clock), .CLR(n2173), .Q(
        reg0[4]) );
  fdef2a6 \reg0_reg[6]  ( .D(N5666), .E(N7156), .CLK(clock), .CLR(n2171), .Q(
        reg0[6]) );
  fdef2a6 \reg0_reg[8]  ( .D(N5670), .E(N7156), .CLK(clock), .CLR(n2169), .Q(
        reg0[8]) );
  fdef2a6 \reg0_reg[10]  ( .D(N5674), .E(N7156), .CLK(clock), .CLR(n2167), .Q(
        reg0[10]) );
  fdef2a6 \reg0_reg[12]  ( .D(N5678), .E(N7156), .CLK(clock), .CLR(n2165), .Q(
        reg0[12]) );
  fdef2a6 \reg0_reg[14]  ( .D(N5682), .E(N7156), .CLK(clock), .CLR(n2163), .Q(
        reg0[14]) );
  fdef2a6 \reg0_reg[16]  ( .D(N5686), .E(N7156), .CLK(clock), .CLR(n2161), .Q(
        reg0[16]) );
  fdef2a6 \reg0_reg[18]  ( .D(N5690), .E(N7156), .CLK(clock), .CLR(n2159), .Q(
        reg0[18]) );
  fdef2a6 \reg0_reg[20]  ( .D(N5694), .E(N7156), .CLK(clock), .CLR(n2157), .Q(
        reg0[20]) );
  fdef2a6 \reg0_reg[22]  ( .D(N5698), .E(N7156), .CLK(clock), .CLR(n2155), .Q(
        reg0[22]) );
  fdef2a6 \reg0_reg[24]  ( .D(N5702), .E(N7156), .CLK(clock), .CLR(n2153), .Q(
        reg0[24]) );
  fdef2a6 \reg0_reg[26]  ( .D(N5706), .E(N7156), .CLK(clock), .CLR(n2151), .Q(
        reg0[26]) );
  fdef2a6 \reg0_reg[28]  ( .D(N5710), .E(N7156), .CLK(clock), .CLR(n2149), .Q(
        reg0[28]) );
  fdef2a6 \reg1_reg[29]  ( .D(N5712), .E(N7188), .CLK(clock), .CLR(n2146), .Q(
        reg1[29]) );
  fdef2a6 \reg1_reg[27]  ( .D(N5708), .E(N7188), .CLK(clock), .CLR(n2150), .Q(
        reg1[27]) );
  fdef2a6 \reg1_reg[25]  ( .D(N5704), .E(N7188), .CLK(clock), .CLR(n2152), .Q(
        reg1[25]) );
  fdef2a6 \reg1_reg[23]  ( .D(N5700), .E(N7188), .CLK(clock), .CLR(n2154), .Q(
        reg1[23]) );
  fdef2a6 \reg1_reg[21]  ( .D(N5696), .E(N7188), .CLK(clock), .CLR(n2156), .Q(
        reg1[21]) );
  fdef2a6 \reg1_reg[20]  ( .D(N5694), .E(N7188), .CLK(clock), .CLR(n2157), .Q(
        reg1[20]) );
  fdef2a6 \reg1_reg[22]  ( .D(N5698), .E(N7188), .CLK(clock), .CLR(n2155), .Q(
        reg1[22]) );
  fdef2a6 \reg1_reg[24]  ( .D(N5702), .E(N7188), .CLK(clock), .CLR(n2153), .Q(
        reg1[24]) );
  fdef2a6 \reg1_reg[26]  ( .D(N5706), .E(N7188), .CLK(clock), .CLR(n2151), .Q(
        reg1[26]) );
  fdef2a6 \reg1_reg[28]  ( .D(N5710), .E(N7188), .CLK(clock), .CLR(n2149), .Q(
        reg1[28]) );
  fdef2a3 \reg1_reg[30]  ( .D(N5778), .E(N7188), .CLK(clock), .CLR(n2147), .Q(
        reg1[30]) );
  fdef2a6 \reg0_reg[30]  ( .D(N5778), .E(N7156), .CLK(clock), .CLR(n2147), .Q(
        reg0[30]) );
  fdef2a6 \reg0_reg[0]  ( .D(N5654), .E(N7156), .CLK(clock), .CLR(n2176), .Q(
        reg0[0]) );
  fdef2a6 \reg2_reg[30]  ( .D(N5778), .E(N7220), .CLK(clock), .CLR(n2147), .Q(
        reg2[30]) );
  fdef2a3 \reg2_reg[31]  ( .D(N5780), .E(N7220), .CLK(clock), .CLR(n2148), .Q(
        reg2[31]) );
  fdef2a6 \reg1_reg[31]  ( .D(N5780), .E(N7188), .CLK(clock), .CLR(n2148), .Q(
        reg1[31]) );
  fdef2a6 \reg0_reg[31]  ( .D(N5780), .E(N7156), .CLK(clock), .CLR(n2147), .Q(
        reg0[31]) );
  fdef2a6 \IR_reg[30]  ( .D(N7055), .E(N7056), .CLK(clock), .CLR(n2178), .Q(
        IR[30]) );
  fdef2a6 \IR_reg[1]  ( .D(N6997), .E(N7056), .CLK(clock), .CLR(n2184), .Q(
        IR[1]) );
  fdef2a6 \IR_reg[2]  ( .D(N6999), .E(N7056), .CLK(clock), .CLR(n2184), .Q(
        IR[2]) );
  fdef2a6 \IR_reg[3]  ( .D(N7001), .E(N7056), .CLK(clock), .CLR(n2183), .Q(
        IR[3]) );
  fdef2a6 \IR_reg[4]  ( .D(N7003), .E(N7056), .CLK(clock), .CLR(n2183), .Q(
        IR[4]) );
  fdef2a6 \IR_reg[8]  ( .D(N7011), .E(N7056), .CLK(clock), .CLR(n2182), .Q(
        IR[8]) );
  fdef2a6 \IR_reg[9]  ( .D(N7013), .E(N7056), .CLK(clock), .CLR(n2182), .Q(
        IR[9]) );
  fdef2a6 \IR_reg[22]  ( .D(N7039), .E(N7056), .CLK(clock), .CLR(n2180), .Q(
        IR[22]) );
  fdef2a6 \IR_reg[23]  ( .D(N7041), .E(N7056), .CLK(clock), .CLR(n2179), .Q(
        IR[23]) );
  fdef2a6 \IR_reg[24]  ( .D(N7043), .E(N7056), .CLK(clock), .CLR(n2179), .Q(
        IR[24]) );
  fdef2a6 \IR_reg[26]  ( .D(N7047), .E(N7056), .CLK(clock), .CLR(n2179), .Q(
        IR[26]) );
  fdef2a6 \IR_reg[27]  ( .D(N7049), .E(N7056), .CLK(clock), .CLR(n2179), .Q(
        IR[27]) );
  fdef2a6 \IR_reg[28]  ( .D(N7051), .E(N7056), .CLK(clock), .CLR(n2178), .Q(
        IR[28]) );
  fdef2a6 \IR_reg[29]  ( .D(N7053), .E(N7056), .CLK(clock), .CLR(n2178), .Q(
        IR[29]) );
  fdef2a6 \IR_reg[5]  ( .D(N7005), .E(N7056), .CLK(clock), .CLR(n2183), .Q(
        IR[5]) );
  fdef2a6 \IR_reg[6]  ( .D(N7007), .E(N7056), .CLK(clock), .CLR(n2183), .Q(
        IR[6]) );
  fdef2a6 \IR_reg[7]  ( .D(N7009), .E(N7056), .CLK(clock), .CLR(n2183), .Q(
        IR[7]) );
  fdef2a6 \IR_reg[10]  ( .D(N7015), .E(N7056), .CLK(clock), .CLR(n2182), .Q(
        IR[10]) );
  fdef2a6 \IR_reg[11]  ( .D(N7017), .E(N7056), .CLK(clock), .CLR(n2182), .Q(
        IR[11]) );
  fdef2a6 \IR_reg[12]  ( .D(N7019), .E(N7056), .CLK(clock), .CLR(n2182), .Q(
        IR[12]) );
  fdef2a6 \IR_reg[13]  ( .D(N7021), .E(N7056), .CLK(clock), .CLR(n2181), .Q(
        IR[13]) );
  fdef2a6 \IR_reg[14]  ( .D(N7023), .E(N7056), .CLK(clock), .CLR(n2181), .Q(
        IR[14]) );
  fdef2a6 \IR_reg[15]  ( .D(N7025), .E(N7056), .CLK(clock), .CLR(n2181), .Q(
        IR[15]) );
  fdef2a6 \IR_reg[16]  ( .D(N7027), .E(N7056), .CLK(clock), .CLR(n2181), .Q(
        IR[16]) );
  fdef2a6 \IR_reg[17]  ( .D(N7029), .E(N7056), .CLK(clock), .CLR(n2181), .Q(
        IR[17]) );
  fdef2a6 \IR_reg[18]  ( .D(N7031), .E(N7056), .CLK(clock), .CLR(n2180), .Q(
        IR[18]) );
  fdef2a6 \IR_reg[19]  ( .D(N7033), .E(N7056), .CLK(clock), .CLR(n2180), .Q(
        IR[19]) );
  fdef2a6 \IR_reg[20]  ( .D(N7035), .E(N7056), .CLK(clock), .CLR(n2180), .Q(
        IR[20]) );
  fdef2a6 \IR_reg[21]  ( .D(N7037), .E(N7056), .CLK(clock), .CLR(n2180), .Q(
        IR[21]) );
  fdef2a6 \IR_reg[25]  ( .D(N7045), .E(N7056), .CLK(clock), .CLR(n2179), .Q(
        IR[25]) );
  fdef2a6 \reg3_reg[28]  ( .D(N6920), .E(state), .CLK(clock), .CLR(n2148), .Q(
        reg3[28]) );
  fdef2a6 \reg3_reg[20]  ( .D(N6912), .E(state), .CLK(clock), .CLR(n2156), .Q(
        reg3[20]) );
  fdef2a6 \reg3_reg[21]  ( .D(N6913), .E(state), .CLK(clock), .CLR(n2155), .Q(
        reg3[21]) );
  fdef2a6 \reg3_reg[22]  ( .D(N6914), .E(state), .CLK(clock), .CLR(n2154), .Q(
        reg3[22]) );
  fdef2a6 \reg3_reg[23]  ( .D(N6915), .E(state), .CLK(clock), .CLR(n2153), .Q(
        reg3[23]) );
  fdef2a6 \reg3_reg[24]  ( .D(N6916), .E(state), .CLK(clock), .CLR(n2152), .Q(
        reg3[24]) );
  fdef2a6 \reg3_reg[25]  ( .D(N6917), .E(state), .CLK(clock), .CLR(n2151), .Q(
        reg3[25]) );
  fdef2a6 \reg3_reg[26]  ( .D(N6918), .E(state), .CLK(clock), .CLR(n2150), .Q(
        reg3[26]) );
  fdef2a6 \reg3_reg[27]  ( .D(N6919), .E(state), .CLK(clock), .CLR(n2149), .Q(
        reg3[27]) );
  fdef2a6 B_reg ( .D(N6754), .E(N7124), .CLK(clock), .CLR(n2177), .Q(B) );
  fdef2a6 \reg3_reg[4]  ( .D(N6896), .E(state), .CLK(clock), .CLR(n2172), .Q(
        reg3[4]) );
  fdef2a6 \reg3_reg[5]  ( .D(N6897), .E(state), .CLK(clock), .CLR(n2171), .Q(
        reg3[5]) );
  fdef2a6 \reg3_reg[6]  ( .D(N6898), .E(state), .CLK(clock), .CLR(n2170), .Q(
        reg3[6]) );
  fdef2a6 \reg3_reg[7]  ( .D(N6899), .E(state), .CLK(clock), .CLR(n2169), .Q(
        reg3[7]) );
  fdef2a6 \reg3_reg[8]  ( .D(N6900), .E(state), .CLK(clock), .CLR(n2168), .Q(
        reg3[8]) );
  fdef2a6 \reg3_reg[9]  ( .D(N6901), .E(state), .CLK(clock), .CLR(n2167), .Q(
        reg3[9]) );
  fdef2a6 \reg3_reg[10]  ( .D(N6902), .E(state), .CLK(clock), .CLR(n2166), .Q(
        reg3[10]) );
  fdef2a6 \reg3_reg[11]  ( .D(N6903), .E(state), .CLK(clock), .CLR(n2165), .Q(
        reg3[11]) );
  fdef2a6 \reg3_reg[12]  ( .D(N6904), .E(state), .CLK(clock), .CLR(n2164), .Q(
        reg3[12]) );
  fdef2a6 \reg3_reg[13]  ( .D(N6905), .E(state), .CLK(clock), .CLR(n2163), .Q(
        reg3[13]) );
  fdef2a6 \reg3_reg[14]  ( .D(N6906), .E(state), .CLK(clock), .CLR(n2162), .Q(
        reg3[14]) );
  fdef2a6 \reg3_reg[15]  ( .D(N6907), .E(state), .CLK(clock), .CLR(n2161), .Q(
        reg3[15]) );
  fdef2a6 \reg3_reg[16]  ( .D(N6908), .E(state), .CLK(clock), .CLR(n2160), .Q(
        reg3[16]) );
  fdef2a6 \reg3_reg[17]  ( .D(N6909), .E(state), .CLK(clock), .CLR(n2159), .Q(
        reg3[17]) );
  fdef2a6 \reg3_reg[18]  ( .D(N6910), .E(state), .CLK(clock), .CLR(n2158), .Q(
        reg3[18]) );
  fdef2a6 \reg3_reg[19]  ( .D(N6911), .E(state), .CLK(clock), .CLR(n2157), .Q(
        reg3[19]) );
  fdef2a6 \IR_reg[0]  ( .D(N6995), .E(N7056), .CLK(clock), .CLR(n2184), .Q(
        IR[0]) );
  fdef2a6 \reg3_reg[1]  ( .D(N6893), .E(state), .CLK(clock), .CLR(n2175), .Q(
        reg3[1]) );
  fdef2a6 \reg3_reg[2]  ( .D(N6894), .E(state), .CLK(clock), .CLR(n2174), .Q(
        reg3[2]) );
  fdef2a6 \reg3_reg[0]  ( .D(N6892), .E(state), .CLK(clock), .CLR(n2176), .Q(
        reg3[0]) );
  fdef2a6 \reg3_reg[3]  ( .D(N6895), .E(state), .CLK(clock), .CLR(n2173), .Q(
        reg3[3]) );
  fdef2a6 \reg1_reg[17]  ( .D(N5688), .E(N7188), .CLK(clock), .CLR(n2160), .Q(
        reg1[17]) );
  fdef2a6 \reg1_reg[15]  ( .D(N5684), .E(N7188), .CLK(clock), .CLR(n2162), .Q(
        reg1[15]) );
  fdef2a6 \reg1_reg[13]  ( .D(N5680), .E(N7188), .CLK(clock), .CLR(n2164), .Q(
        reg1[13]) );
  fdef2a6 \reg1_reg[11]  ( .D(N5676), .E(N7188), .CLK(clock), .CLR(n2166), .Q(
        reg1[11]) );
  fdef2a6 \reg1_reg[3]  ( .D(N5660), .E(N7188), .CLK(clock), .CLR(n2174), .Q(
        reg1[3]) );
  fdef2a6 \reg1_reg[1]  ( .D(N5656), .E(N7188), .CLK(clock), .CLR(n2176), .Q(
        reg1[1]) );
  fdef2a6 \reg1_reg[2]  ( .D(N5658), .E(N7188), .CLK(clock), .CLR(n2175), .Q(
        reg1[2]) );
  fdef2a6 \reg1_reg[10]  ( .D(N5674), .E(N7188), .CLK(clock), .CLR(n2167), .Q(
        reg1[10]) );
  fdef2a6 \reg1_reg[12]  ( .D(N5678), .E(N7188), .CLK(clock), .CLR(n2165), .Q(
        reg1[12]) );
  fdef2a6 \reg1_reg[14]  ( .D(N5682), .E(N7188), .CLK(clock), .CLR(n2163), .Q(
        reg1[14]) );
  fdef2a6 \reg1_reg[16]  ( .D(N5686), .E(N7188), .CLK(clock), .CLR(n2161), .Q(
        reg1[16]) );
  fdef2a6 \reg1_reg[18]  ( .D(N5690), .E(N7188), .CLK(clock), .CLR(n2159), .Q(
        reg1[18]) );
  fdef2a6 \reg1_reg[9]  ( .D(N5672), .E(N7188), .CLK(clock), .CLR(n2168), .Q(
        reg1[9]) );
  fdef2a6 \reg1_reg[7]  ( .D(N5668), .E(N7188), .CLK(clock), .CLR(n2170), .Q(
        reg1[7]) );
  fdef2a6 \reg1_reg[5]  ( .D(N5664), .E(N7188), .CLK(clock), .CLR(n2172), .Q(
        reg1[5]) );
  fdef2a6 \reg1_reg[4]  ( .D(N5662), .E(N7188), .CLK(clock), .CLR(n2173), .Q(
        reg1[4]) );
  fdef2a6 \reg1_reg[6]  ( .D(N5666), .E(N7188), .CLK(clock), .CLR(n2171), .Q(
        reg1[6]) );
  fdef2a6 \reg1_reg[8]  ( .D(N5670), .E(N7188), .CLK(clock), .CLR(n2169), .Q(
        reg1[8]) );
  fdef2a6 \reg2_reg[1]  ( .D(N5720), .E(N7220), .CLK(clock), .CLR(n2175), .Q(
        reg2[1]) );
  fdef2a6 \reg2_reg[2]  ( .D(N5722), .E(N7220), .CLK(clock), .CLR(n2174), .Q(
        reg2[2]) );
  fdef2a6 \reg2_reg[3]  ( .D(N5724), .E(N7220), .CLK(clock), .CLR(n2173), .Q(
        reg2[3]) );
  fdef2a6 \reg2_reg[10]  ( .D(N5738), .E(N7220), .CLK(clock), .CLR(n2166), .Q(
        reg2[10]) );
  fdef2a6 \reg2_reg[11]  ( .D(N5740), .E(N7220), .CLK(clock), .CLR(n2165), .Q(
        reg2[11]) );
  fdef2a6 \reg2_reg[12]  ( .D(N5742), .E(N7220), .CLK(clock), .CLR(n2164), .Q(
        reg2[12]) );
  fdef2a6 \reg2_reg[13]  ( .D(N5744), .E(N7220), .CLK(clock), .CLR(n2163), .Q(
        reg2[13]) );
  fdef2a6 \reg2_reg[14]  ( .D(N5746), .E(N7220), .CLK(clock), .CLR(n2162), .Q(
        reg2[14]) );
  fdef2a6 \reg2_reg[15]  ( .D(N5748), .E(N7220), .CLK(clock), .CLR(n2161), .Q(
        reg2[15]) );
  fdef2a6 \reg2_reg[16]  ( .D(N5750), .E(N7220), .CLK(clock), .CLR(n2160), .Q(
        reg2[16]) );
  fdef2a6 \reg2_reg[17]  ( .D(N5752), .E(N7220), .CLK(clock), .CLR(n2159), .Q(
        reg2[17]) );
  fdef2a6 \reg2_reg[18]  ( .D(N5754), .E(N7220), .CLK(clock), .CLR(n2158), .Q(
        reg2[18]) );
  fdef2a6 \reg2_reg[19]  ( .D(N5756), .E(N7220), .CLK(clock), .CLR(n2157), .Q(
        reg2[19]) );
  fdef2a6 \reg1_reg[19]  ( .D(N5692), .E(N7188), .CLK(clock), .CLR(n2158), .Q(
        reg1[19]) );
  fdef2a6 \reg2_reg[4]  ( .D(N5726), .E(N7220), .CLK(clock), .CLR(n2172), .Q(
        reg2[4]) );
  fdef2a6 \reg2_reg[5]  ( .D(N5728), .E(N7220), .CLK(clock), .CLR(n2171), .Q(
        reg2[5]) );
  fdef2a6 \reg2_reg[6]  ( .D(N5730), .E(N7220), .CLK(clock), .CLR(n2170), .Q(
        reg2[6]) );
  fdef2a6 \reg2_reg[7]  ( .D(N5732), .E(N7220), .CLK(clock), .CLR(n2169), .Q(
        reg2[7]) );
  fdef2a6 \reg2_reg[8]  ( .D(N5734), .E(N7220), .CLK(clock), .CLR(n2168), .Q(
        reg2[8]) );
  fdef2a6 \reg2_reg[9]  ( .D(N5736), .E(N7220), .CLK(clock), .CLR(n2167), .Q(
        reg2[9]) );
  fdef2a6 \reg2_reg[0]  ( .D(N5718), .E(N7220), .CLK(clock), .CLR(n2177), .Q(
        reg2[0]) );
  fdef2a6 \reg1_reg[0]  ( .D(N5654), .E(N7188), .CLK(clock), .CLR(n2177), .Q(
        reg1[0]) );
  fdef2a6 \IR_reg[31]  ( .D(N7057), .E(N7056), .CLK(clock), .CLR(n2184), .Q(
        N325) );
  fdef2a9 state_reg ( .D(N7058), .E(1), .CLK(clock), .CLR(n2184), .Q(state)
         );
  fdef2a3 wr_reg ( .D(N7091), .E(1), .CLK(clock), .CLR(n2178), .Q(wr) );
  fdef2a3 \datao_reg[0]  ( .D(N654), .E(N7091), .CLK(clock), .CLR(n2176), .Q(
        datao[0]) );
  fdef2a3 \datao_reg[1]  ( .D(N655), .E(N7091), .CLK(clock), .CLR(n2175), .Q(
        datao[1]) );
  fdef2a3 \datao_reg[2]  ( .D(N656), .E(N7091), .CLK(clock), .CLR(n2174), .Q(
        datao[2]) );
  fdef2a3 \datao_reg[3]  ( .D(N657), .E(N7091), .CLK(clock), .CLR(n2173), .Q(
        datao[3]) );
  fdef2a3 \datao_reg[4]  ( .D(N658), .E(N7091), .CLK(clock), .CLR(n2172), .Q(
        datao[4]) );
  fdef2a3 \datao_reg[5]  ( .D(N659), .E(N7091), .CLK(clock), .CLR(n2171), .Q(
        datao[5]) );
  fdef2a3 \datao_reg[6]  ( .D(N660), .E(N7091), .CLK(clock), .CLR(n2170), .Q(
        datao[6]) );
  fdef2a3 \datao_reg[7]  ( .D(N661), .E(N7091), .CLK(clock), .CLR(n2169), .Q(
        datao[7]) );
  fdef2a3 \datao_reg[8]  ( .D(N662), .E(N7091), .CLK(clock), .CLR(n2168), .Q(
        datao[8]) );
  fdef2a3 \datao_reg[9]  ( .D(N663), .E(N7091), .CLK(clock), .CLR(n2167), .Q(
        datao[9]) );
  fdef2a3 \datao_reg[10]  ( .D(N664), .E(N7091), .CLK(clock), .CLR(n2166), .Q(
        datao[10]) );
  fdef2a3 \datao_reg[11]  ( .D(N665), .E(N7091), .CLK(clock), .CLR(n2165), .Q(
        datao[11]) );
  fdef2a3 \datao_reg[12]  ( .D(N666), .E(N7091), .CLK(clock), .CLR(n2164), .Q(
        datao[12]) );
  fdef2a3 \datao_reg[13]  ( .D(N667), .E(N7091), .CLK(clock), .CLR(n2163), .Q(
        datao[13]) );
  fdef2a3 \datao_reg[14]  ( .D(N668), .E(N7091), .CLK(clock), .CLR(n2162), .Q(
        datao[14]) );
  fdef2a3 \datao_reg[15]  ( .D(N669), .E(N7091), .CLK(clock), .CLR(n2161), .Q(
        datao[15]) );
  fdef2a3 \datao_reg[16]  ( .D(N670), .E(N7091), .CLK(clock), .CLR(n2160), .Q(
        datao[16]) );
  fdef2a3 \datao_reg[17]  ( .D(N671), .E(N7091), .CLK(clock), .CLR(n2159), .Q(
        datao[17]) );
  fdef2a3 \datao_reg[18]  ( .D(N672), .E(N7091), .CLK(clock), .CLR(n2158), .Q(
        datao[18]) );
  fdef2a3 \datao_reg[19]  ( .D(N673), .E(N7091), .CLK(clock), .CLR(n2157), .Q(
        datao[19]) );
  fdef2a3 \datao_reg[20]  ( .D(N674), .E(N7091), .CLK(clock), .CLR(n2156), .Q(
        datao[20]) );
  fdef2a3 \datao_reg[21]  ( .D(N675), .E(N7091), .CLK(clock), .CLR(n2155), .Q(
        datao[21]) );
  fdef2a3 \datao_reg[22]  ( .D(N676), .E(N7091), .CLK(clock), .CLR(n2154), .Q(
        datao[22]) );
  fdef2a3 \datao_reg[23]  ( .D(N677), .E(N7091), .CLK(clock), .CLR(n2153), .Q(
        datao[23]) );
  fdef2a3 \datao_reg[24]  ( .D(N678), .E(N7091), .CLK(clock), .CLR(n2152), .Q(
        datao[24]) );
  fdef2a3 \datao_reg[25]  ( .D(N679), .E(N7091), .CLK(clock), .CLR(n2151), .Q(
        datao[25]) );
  fdef2a3 \datao_reg[26]  ( .D(N680), .E(N7091), .CLK(clock), .CLR(n2150), .Q(
        datao[26]) );
  fdef2a3 \datao_reg[27]  ( .D(N681), .E(N7091), .CLK(clock), .CLR(n2149), .Q(
        datao[27]) );
  fdef2a3 \datao_reg[28]  ( .D(N682), .E(N7091), .CLK(clock), .CLR(n2148), .Q(
        datao[28]) );
  fdef2a6 \datao_reg[29]  ( .D(N683), .E(N7091), .CLK(clock), .CLR(n2146), .Q(
        datao[29]) );
  fdef2a3 \datao_reg[30]  ( .D(N684), .E(N7091), .CLK(clock), .CLR(n2146), .Q(
        datao[30]) );
  fdef2a3 \datao_reg[31]  ( .D(N685), .E(N7091), .CLK(clock), .CLR(n2147), .Q(
        datao[31]) );
  fdef2a6 \addr_reg[19]  ( .D(N6992), .E(N6991), .CLK(clock), .CLR(n2204), .Q(
        addr[19]) );
  fdef2a6 \addr_reg[17]  ( .D(N6988), .E(N6991), .CLK(clock), .CLR(n2203), .Q(
        addr[17]) );
  fdef2a6 \addr_reg[15]  ( .D(N6984), .E(N6991), .CLK(clock), .CLR(n2205), .Q(
        addr[15]) );
  fdef2a6 \addr_reg[13]  ( .D(N6980), .E(N6991), .CLK(clock), .CLR(n2143), .Q(
        addr[13]) );
  fdef2a6 \addr_reg[11]  ( .D(N6976), .E(N6991), .CLK(clock), .CLR(n2143), .Q(
        addr[11]) );
  fdef2a6 \addr_reg[9]  ( .D(N6972), .E(N6991), .CLK(clock), .CLR(n2144), .Q(
        addr[9]) );
  fdef2a6 \addr_reg[7]  ( .D(N6968), .E(N6991), .CLK(clock), .CLR(n2144), .Q(
        addr[7]) );
  fdef2a6 \addr_reg[5]  ( .D(N6964), .E(N6991), .CLK(clock), .CLR(n2144), .Q(
        addr[5]) );
  fdef2a6 \addr_reg[3]  ( .D(N6960), .E(N6991), .CLK(clock), .CLR(n2145), .Q(
        addr[3]) );
  fdef2a6 \addr_reg[1]  ( .D(N6956), .E(N6991), .CLK(clock), .CLR(n2145), .Q(
        addr[1]) );
  fdef2a6 \addr_reg[0]  ( .D(N6954), .E(N6991), .CLK(clock), .CLR(n2145), .Q(
        addr[0]) );
  fdef2a6 \addr_reg[2]  ( .D(N6958), .E(N6991), .CLK(clock), .CLR(n2145), .Q(
        addr[2]) );
  fdef2a6 \addr_reg[4]  ( .D(N6962), .E(N6991), .CLK(clock), .CLR(n2145), .Q(
        addr[4]) );
  fdef2a6 \addr_reg[6]  ( .D(N6966), .E(N6991), .CLK(clock), .CLR(n2144), .Q(
        addr[6]) );
  fdef2a6 \addr_reg[8]  ( .D(N6970), .E(N6991), .CLK(clock), .CLR(n2144), .Q(
        addr[8]) );
  fdef2a6 \addr_reg[10]  ( .D(N6974), .E(N6991), .CLK(clock), .CLR(n2143), .Q(
        addr[10]) );
  fdef2a6 \addr_reg[12]  ( .D(N6978), .E(N6991), .CLK(clock), .CLR(n2143), .Q(
        addr[12]) );
  fdef2a6 \addr_reg[14]  ( .D(N6982), .E(N6991), .CLK(clock), .CLR(n2143), .Q(
        addr[14]) );
  fdef2a6 \addr_reg[16]  ( .D(N6986), .E(N6991), .CLK(clock), .CLR(n2199), .Q(
        addr[16]) );
  fdef2a6 \addr_reg[18]  ( .D(N6990), .E(N6991), .CLK(clock), .CLR(n425), .Q(
        addr[18]) );
  fdef2a6 rd_reg ( .D(N6993), .E(1), .CLK(clock), .CLR(n2178), .Q(rd) );
  and2a3 U2231 ( .A(N548), .B(n2234), .Y(n2239) );
  and2a3 U2232 ( .A(N550), .B(n2234), .Y(n2245) );
  and2a3 U2233 ( .A(n3041), .B(n3053), .Y(n3046) );
  and2a3 U2234 ( .A(n2622), .B(N537), .Y(n2629) );
  and2a3 U2235 ( .A(n2622), .B(N553), .Y(n2746) );
  and2a3 U2236 ( .A(n2622), .B(N555), .Y(n2764) );
  and2a3 U2237 ( .A(n2622), .B(N554), .Y(n2757) );
  and2a3 U2238 ( .A(n2595), .B(N941), .Y(\U3/U1/Z_2 ) );
  and2a3 U2239 ( .A(n2595), .B(N958), .Y(\U3/U1/Z_19 ) );
  and2a3 U2240 ( .A(n2595), .B(N957), .Y(\U3/U1/Z_18 ) );
  and2a3 U2241 ( .A(n2595), .B(N956), .Y(\U3/U1/Z_17 ) );
  and2a3 U2242 ( .A(n2595), .B(N955), .Y(\U3/U1/Z_16 ) );
  and2a3 U2243 ( .A(n2595), .B(N953), .Y(\U3/U1/Z_14 ) );
  and2a3 U2244 ( .A(n2595), .B(N952), .Y(\U3/U1/Z_13 ) );
  and2a3 U2245 ( .A(n2595), .B(N951), .Y(\U3/U1/Z_12 ) );
  and2a3 U2246 ( .A(n2595), .B(N949), .Y(\U3/U1/Z_10 ) );
  and2a3 U2247 ( .A(n2595), .B(N948), .Y(\U3/U1/Z_9 ) );
  and2a3 U2248 ( .A(n2595), .B(N947), .Y(\U3/U1/Z_8 ) );
  and2a3 U2249 ( .A(n2595), .B(N945), .Y(\U3/U1/Z_6 ) );
  and2a3 U2250 ( .A(n2595), .B(N944), .Y(\U3/U1/Z_5 ) );
  and2a3 U2251 ( .A(n2595), .B(N943), .Y(\U3/U1/Z_4 ) );
  and2a3 U2252 ( .A(n2622), .B(N543), .Y(n2671) );
  mx2a3 U2253 ( .D0(N305), .D1(IR[12]), .S(n3731), .Y(N543) );
  and2a3 U2254 ( .A(n2622), .B(N542), .Y(n2664) );
  mx2a3 U2255 ( .D0(N306), .D1(IR[13]), .S(n3731), .Y(N542) );
  mx2a3 U2256 ( .D0(N307), .D1(IR[14]), .S(n3731), .Y(N541) );
  and2a3 U2257 ( .A(N552), .B(n2234), .Y(n2252) );
  mx2a3 U2258 ( .D0(IR[3]), .D1(N296), .S(N325), .Y(N552) );
  mx2a3 U2259 ( .D0(N304), .D1(IR[11]), .S(n3731), .Y(N544) );
  inv1a3 U2260 ( .A(N678), .Y(n2265) );
  xor2a6 U2261 ( .A(n3023), .B(n3024), .Y(n2605) );
  and2a3 U2262 ( .A(N547), .B(n2234), .Y(n2236) );
  mx2a3 U2263 ( .D0(IR[8]), .D1(N301), .S(N325), .Y(N547) );
  and2a3 U2264 ( .A(n2622), .B(N538), .Y(n2636) );
  mx2a3 U2265 ( .D0(N310), .D1(IR[17]), .S(n3731), .Y(N538) );
  inv1a3 U2266 ( .A(N679), .Y(n2263) );
  and2a3 U2267 ( .A(N551), .B(n2234), .Y(n2248) );
  mx2a3 U2268 ( .D0(IR[4]), .D1(N297), .S(N325), .Y(N551) );
  mx2a3 U2269 ( .D0(N308), .D1(IR[15]), .S(n3731), .Y(N540) );
  inv1a3 U2270 ( .A(n2849), .Y(n2792) );
  inv1a3 U2271 ( .A(N674), .Y(n2273) );
  inv1a3 U2272 ( .A(N676), .Y(n2269) );
  inv1a3 U2273 ( .A(N680), .Y(n2261) );
  inv1a3 U2274 ( .A(N675), .Y(n2271) );
  inv1a3 U2275 ( .A(N677), .Y(n2267) );
  inv1a3 U2276 ( .A(N681), .Y(n2259) );
  inv1a3 U2277 ( .A(N673), .Y(n2278) );
  and2a3 U2278 ( .A(n3043), .B(n3002), .Y(n3049) );
  and2a3 U2279 ( .A(n3002), .B(n3046), .Y(n3036) );
  xor2a6 U2280 ( .A(n3728), .B(n3737), .Y(n3002) );
  and2a3 U2281 ( .A(n2622), .B(N546), .Y(n2692) );
  and2a3 U2282 ( .A(N546), .B(n2234), .Y(n2232) );
  mx2a3 U2283 ( .D0(IR[9]), .D1(N302), .S(N325), .Y(N546) );
  and2a3 U2284 ( .A(n2622), .B(N539), .Y(n2643) );
  mx2a3 U2285 ( .D0(N309), .D1(IR[16]), .S(n3731), .Y(N539) );
  and2a6 U2286 ( .A(n2595), .B(n2314), .Y(n2791) );
  oa1f3 U2287 ( .A(n2776), .B(n2777), .C(n2778), .Y(n2622) );
  and2a6 U2288 ( .A(n3113), .B(n3036), .Y(n2998) );
  xor2a6 U2289 ( .A(n3730), .B(n3735), .Y(n3043) );
  or3a2 U2290 ( .A(n3099), .B(n3100), .C(n3101), .Y(N685) );
  mx2a3 U2291 ( .D0(IR[1]), .D1(N294), .S(N325), .Y(N554) );
  mx2a3 U2292 ( .D0(N311), .D1(IR[18]), .S(n3731), .Y(N537) );
  inv1a3 U2293 ( .A(n2555), .Y(n2552) );
  or4a6 U2294 ( .A(n3671), .B(n3672), .C(n3673), .D(n3674), .Y(N655) );
  and2a6 U2295 ( .A(n2314), .B(n2317), .Y(n2230) );
  and3a3 U2296 ( .A(n2771), .B(n2316), .C(n2596), .Y(n2618) );
  and4a6 U2297 ( .A(n3113), .B(n3050), .C(n3053), .D(n3002), .Y(n2580) );
  inv1a2 U2298 ( .A(n3043), .Y(n3053) );
  inv1a3 U2299 ( .A(N682), .Y(n2257) );
  and4a6 U2300 ( .A(n3720), .B(n3004), .C(n3041), .D(n3043), .Y(n3001) );
  inv1a3 U2301 ( .A(n3050), .Y(n3041) );
  inv1a3 U2302 ( .A(n2319), .Y(n2338) );
  or4a6 U2303 ( .A(n3255), .B(n3256), .C(n3257), .D(n3258), .Y(N676) );
  or4a6 U2304 ( .A(n3179), .B(n3180), .C(n3181), .D(n3182), .Y(N680) );
  or4a6 U2305 ( .A(n3236), .B(n3237), .C(n3238), .D(n3239), .Y(N677) );
  or4a6 U2306 ( .A(n3160), .B(n3161), .C(n3162), .D(n3163), .Y(N681) );
  or4a6 U2307 ( .A(n3312), .B(n3313), .C(n3314), .D(n3315), .Y(N673) );
  or4a6 U2308 ( .A(n3293), .B(n3294), .C(n3295), .D(n3296), .Y(N674) );
  or4a6 U2309 ( .A(n3217), .B(n3218), .C(n3219), .D(n3220), .Y(N678) );
  or4a6 U2310 ( .A(n3274), .B(n3275), .C(n3276), .D(n3277), .Y(N675) );
  or4a6 U2311 ( .A(n3198), .B(n3199), .C(n3200), .D(n3201), .Y(N679) );
  or4a6 U2312 ( .A(n3651), .B(n3652), .C(n3653), .D(n3654), .Y(N656) );
  or4a6 U2313 ( .A(n3631), .B(n3632), .C(n3633), .D(n3634), .Y(N657) );
  or4a6 U2314 ( .A(n3571), .B(n3572), .C(n3573), .D(n3574), .Y(N660) );
  or4a6 U2315 ( .A(n3551), .B(n3552), .C(n3553), .D(n3554), .Y(N661) );
  or4a6 U2316 ( .A(n3491), .B(n3492), .C(n3493), .D(n3494), .Y(N664) );
  or4a6 U2317 ( .A(n3471), .B(n3472), .C(n3473), .D(n3474), .Y(N665) );
  or4a6 U2318 ( .A(n3411), .B(n3412), .C(n3413), .D(n3414), .Y(N668) );
  or4a6 U2319 ( .A(n3391), .B(n3392), .C(n3393), .D(n3394), .Y(N669) );
  or4a6 U2320 ( .A(n3331), .B(n3332), .C(n3333), .D(n3334), .Y(N672) );
  mx2a3 U2321 ( .D0(IR[0]), .D1(N293), .S(N325), .Y(N555) );
  or4a6 U2322 ( .A(n3591), .B(n3592), .C(n3593), .D(n3594), .Y(N659) );
  or4a6 U2323 ( .A(n3511), .B(n3512), .C(n3513), .D(n3514), .Y(N663) );
  or4a6 U2324 ( .A(n3431), .B(n3432), .C(n3433), .D(n3434), .Y(N667) );
  or4a6 U2325 ( .A(n3351), .B(n3352), .C(n3353), .D(n3354), .Y(N671) );
  or4a6 U2326 ( .A(n3611), .B(n3612), .C(n3613), .D(n3614), .Y(N658) );
  or4a6 U2327 ( .A(n3451), .B(n3452), .C(n3453), .D(n3454), .Y(N666) );
  or4a6 U2328 ( .A(n3371), .B(n3372), .C(n3373), .D(n3374), .Y(N670) );
  or4a6 U2329 ( .A(n3531), .B(n3532), .C(n3533), .D(n3534), .Y(N662) );
  xor2a6 U2330 ( .A(N536), .B(n3027), .Y(n3050) );
  mx2a3 U2331 ( .D0(N312), .D1(IR[19]), .S(n3731), .Y(N536) );
  or4a6 U2332 ( .A(n3692), .B(n3693), .C(n3694), .D(n3695), .Y(N654) );
  and3a3 U2333 ( .A(n2313), .B(n2772), .C(n2596), .Y(n2620) );
  and3a9 U2334 ( .A(n3720), .B(n3043), .C(n3113), .Y(n2996) );
  and3a9 U2335 ( .A(n2999), .B(n2314), .C(n2583), .Y(n2790) );
  or4a6 U2336 ( .A(n3138), .B(n3139), .C(n3140), .D(n3141), .Y(N682) );
  mx2a3 U2337 ( .D0(IR[2]), .D1(N295), .S(N325), .Y(N553) );
  oa1f2 U2338 ( .A(n2471), .B(reg2[19]), .C(n2496), .Y(n2492) );
  inv1a3 U2339 ( .A(n2395), .Y(N940) );
  inv1a3 U2340 ( .A(n2556), .Y(n2536) );
  and2a6 U2341 ( .A(n2465), .B(n2338), .Y(n2400) );
  and3a3 U2342 ( .A(n2313), .B(n2314), .C(n2315), .Y(n2206) );
  ao1f3 U2343 ( .A(N7058), .B(n2773), .C(n2774), .Y(n2621) );
  ao1f9 U2344 ( .A(n2623), .B(n2592), .C(n2610), .Y(N6991) );
  or3a6 U2345 ( .A(n2992), .B(n2993), .C(n2462), .Y(n2787) );
  and3a9 U2346 ( .A(n3720), .B(n3004), .C(n3046), .Y(n2997) );
  xor2a6 U2347 ( .A(n3729), .B(n3736), .Y(n3004) );
  inv1a2 U2348 ( .A(n3002), .Y(n3720) );
  and3a9 U2349 ( .A(n2599), .B(n2603), .C(n2601), .Y(N7156) );
  and3a9 U2350 ( .A(n3113), .B(n3053), .C(n3056), .Y(n2597) );
  or3a2 U2351 ( .A(n3102), .B(n3103), .C(n3104), .Y(N684) );
  mx2a3 U2352 ( .D0(N298), .D1(IR[5]), .S(n3731), .Y(N550) );
  mx2a3 U2353 ( .D0(N299), .D1(IR[6]), .S(n3731), .Y(N549) );
  mx2a3 U2354 ( .D0(N300), .D1(IR[7]), .S(n3731), .Y(N548) );
  mx2a3 U2355 ( .D0(N303), .D1(IR[10]), .S(n3731), .Y(N545) );
  inv1a3 U2356 ( .A(N325), .Y(n3731) );
  and3a3 U2357 ( .A(n2771), .B(n2315), .C(n2596), .Y(n2619) );
  and3a3 U2358 ( .A(n2313), .B(n2314), .C(n2316), .Y(n2208) );
  and2a6 U2359 ( .A(n3699), .B(n3697), .Y(n3095) );
  and2a6 U2360 ( .A(n3698), .B(n3696), .Y(n3097) );
  ao1f3 U2361 ( .A(n2463), .B(n2585), .C(n2587), .Y(n2471) );
  inv1a6 U2362 ( .A(n2579), .Y(n2539) );
  or2a6 U2363 ( .A(n3691), .B(n2464), .Y(n3137) );
  inv1a6 U2364 ( .A(n2322), .Y(n2401) );
  ao1f6 U2365 ( .A(n2590), .B(n2591), .C(n2592), .Y(n2319) );
  ao1a6 U2366 ( .A(n3006), .B(n2583), .C(\U3/U2/Z_0 ), .Y(n2595) );
  and3a9 U2367 ( .A(n3053), .B(n3004), .C(n3056), .Y(n2582) );
  and3a9 U2368 ( .A(n2602), .B(n2603), .C(n2601), .Y(N7188) );
  and3a9 U2369 ( .A(n3113), .B(n3050), .C(n3049), .Y(n2593) );
  and3a9 U2370 ( .A(n2314), .B(n2755), .C(n2986), .Y(n2789) );
  xor2a6 U2371 ( .A(n3706), .B(n3723), .Y(n2755) );
  inv1a3 U2372 ( .A(n2472), .Y(n2491) );
  or2a6 U2373 ( .A(\U3/U5/Z_0 ), .B(n2530), .Y(n2472) );
  inv1a3 U2374 ( .A(n2365), .Y(N958) );
  inv1a3 U2375 ( .A(n2371), .Y(N956) );
  inv1a3 U2376 ( .A(n2383), .Y(N952) );
  inv1a3 U2377 ( .A(n2318), .Y(N948) );
  inv1a3 U2378 ( .A(n2332), .Y(N944) );
  inv1a3 U2379 ( .A(n2335), .Y(N943) );
  inv1a3 U2380 ( .A(n2323), .Y(N947) );
  inv1a3 U2381 ( .A(n2386), .Y(N951) );
  inv1a3 U2382 ( .A(n2374), .Y(N955) );
  inv1a3 U2383 ( .A(n2377), .Y(N954) );
  inv1a3 U2384 ( .A(n2389), .Y(N950) );
  inv1a3 U2385 ( .A(n2326), .Y(N946) );
  inv1a3 U2386 ( .A(n2339), .Y(N942) );
  inv1a3 U2387 ( .A(n2362), .Y(N941) );
  inv1a3 U2388 ( .A(n2329), .Y(N945) );
  inv1a3 U2389 ( .A(n2392), .Y(N949) );
  inv1a3 U2390 ( .A(n2380), .Y(N953) );
  inv1a3 U2391 ( .A(n2368), .Y(N957) );
  and2a6 U2392 ( .A(n3696), .B(n3697), .Y(n3096) );
  or2a6 U2393 ( .A(n2208), .B(n2206), .Y(n2234) );
  ao1f3 U2394 ( .A(n2584), .B(n2585), .C(n2586), .Y(n2470) );
  and2a6 U2395 ( .A(n3698), .B(n3699), .Y(n3098) );
  ao1a6 U2396 ( .A(N555), .B(n3143), .C(n3721), .Y(N939) );
  inv1a6 U2397 ( .A(n2317), .Y(n3159) );
  and3a9 U2398 ( .A(n3005), .B(n2314), .C(n2986), .Y(n2788) );
  or3a6 U2399 ( .A(n2462), .B(n2463), .C(n2464), .Y(n2322) );
  inv1a6 U2400 ( .A(state), .Y(N7058) );
  inv1a6 U2401 ( .A(n3007), .Y(\U3/U2/Z_0 ) );
  ao1a6 U2402 ( .A(n2531), .B(n2532), .C(n2533), .Y(\U3/U5/Z_0 ) );
  and3a9 U2403 ( .A(n3004), .B(n3043), .C(n3056), .Y(n3000) );
  or2a6 U2404 ( .A(N325), .B(N7058), .Y(N7056) );
  ao1a6 U2405 ( .A(n2596), .B(n2597), .C(n2598), .Y(N7220) );
  and3a9 U2406 ( .A(n3113), .B(n3041), .C(n3049), .Y(n2581) );
  and3a9 U2407 ( .A(n3046), .B(n3720), .C(n3113), .Y(n2532) );
  inv1a2 U2408 ( .A(n3004), .Y(n3113) );
  or2a6 U2409 ( .A(n2779), .B(n2772), .Y(n2624) );
  and3a9 U2410 ( .A(state), .B(n2605), .C(n2607), .Y(N7091) );
  inv1a6 U2411 ( .A(\U3/U10/Z_0 ), .Y(n2255) );
  and2a9 U2412 ( .A(n2466), .B(n2338), .Y(\U3/U10/Z_0 ) );
  buf1a3 U2413 ( .A(n2198), .Y(n2145) );
  buf1a3 U2414 ( .A(n2198), .Y(n2144) );
  buf1a3 U2415 ( .A(n2198), .Y(n2143) );
  buf1a3 U2416 ( .A(n2197), .Y(n2147) );
  buf1a3 U2417 ( .A(n2187), .Y(n2177) );
  buf1a3 U2418 ( .A(n2197), .Y(n2146) );
  buf1a3 U2419 ( .A(n2197), .Y(n2148) );
  buf1a3 U2420 ( .A(n2196), .Y(n2149) );
  buf1a3 U2421 ( .A(n2196), .Y(n2150) );
  buf1a3 U2422 ( .A(n2196), .Y(n2151) );
  buf1a3 U2423 ( .A(n2195), .Y(n2152) );
  buf1a3 U2424 ( .A(n2195), .Y(n2153) );
  buf1a3 U2425 ( .A(n2195), .Y(n2154) );
  buf1a3 U2426 ( .A(n2194), .Y(n2155) );
  buf1a3 U2427 ( .A(n2194), .Y(n2156) );
  buf1a3 U2428 ( .A(n2194), .Y(n2157) );
  buf1a3 U2429 ( .A(n2193), .Y(n2158) );
  buf1a3 U2430 ( .A(n2193), .Y(n2159) );
  buf1a3 U2431 ( .A(n2193), .Y(n2160) );
  buf1a3 U2432 ( .A(n2192), .Y(n2161) );
  buf1a3 U2433 ( .A(n2192), .Y(n2162) );
  buf1a3 U2434 ( .A(n2192), .Y(n2163) );
  buf1a3 U2435 ( .A(n2191), .Y(n2164) );
  buf1a3 U2436 ( .A(n2191), .Y(n2165) );
  buf1a3 U2437 ( .A(n2191), .Y(n2166) );
  buf1a3 U2438 ( .A(n2190), .Y(n2167) );
  buf1a3 U2439 ( .A(n2190), .Y(n2168) );
  buf1a3 U2440 ( .A(n2190), .Y(n2169) );
  buf1a3 U2441 ( .A(n2189), .Y(n2170) );
  buf1a3 U2442 ( .A(n2189), .Y(n2171) );
  buf1a3 U2443 ( .A(n2189), .Y(n2172) );
  buf1a3 U2444 ( .A(n2188), .Y(n2173) );
  buf1a3 U2445 ( .A(n2188), .Y(n2174) );
  buf1a3 U2446 ( .A(n2188), .Y(n2175) );
  buf1a3 U2447 ( .A(n2187), .Y(n2176) );
  buf1a3 U2448 ( .A(n2186), .Y(n2179) );
  buf1a3 U2449 ( .A(n2186), .Y(n2180) );
  buf1a3 U2450 ( .A(n2186), .Y(n2181) );
  buf1a3 U2451 ( .A(n2185), .Y(n2182) );
  buf1a3 U2452 ( .A(n2185), .Y(n2183) );
  buf1a3 U2453 ( .A(n2187), .Y(n2178) );
  buf1a3 U2454 ( .A(n2185), .Y(n2184) );
  buf1a3 U2455 ( .A(n2199), .Y(n2198) );
  buf1a3 U2456 ( .A(n2199), .Y(n2197) );
  buf1a3 U2457 ( .A(n2200), .Y(n2196) );
  buf1a3 U2458 ( .A(n2200), .Y(n2195) );
  buf1a3 U2459 ( .A(n2200), .Y(n2194) );
  buf1a3 U2460 ( .A(n2201), .Y(n2193) );
  buf1a3 U2461 ( .A(n2201), .Y(n2192) );
  buf1a3 U2462 ( .A(n2201), .Y(n2191) );
  buf1a3 U2463 ( .A(n2202), .Y(n2190) );
  buf1a3 U2464 ( .A(n2202), .Y(n2189) );
  buf1a3 U2465 ( .A(n2202), .Y(n2188) );
  buf1a3 U2466 ( .A(n2203), .Y(n2186) );
  buf1a3 U2467 ( .A(n2203), .Y(n2187) );
  buf1a3 U2468 ( .A(n2203), .Y(n2185) );
  buf1a3 U2469 ( .A(n2205), .Y(n2199) );
  buf1a3 U2470 ( .A(n2205), .Y(n2200) );
  buf1a3 U2471 ( .A(n2204), .Y(n2201) );
  buf1a3 U2472 ( .A(n2204), .Y(n2202) );
  buf1a3 U2473 ( .A(n2204), .Y(n2203) );
  buf1a3 U2474 ( .A(n425), .Y(n2204) );
  buf1a3 U2475 ( .A(n425), .Y(n2205) );
  inv1a1 U2476 ( .A(reset), .Y(n425) );
  ao1a1 U2477 ( .A(n2206), .B(reg1[9]), .C(n2207), .Y(\U3/U9/Z_9 ) );
  and2a3 U2478 ( .A(n2208), .B(reg2[9]), .Y(n2207) );
  ao1a1 U2479 ( .A(n2206), .B(reg1[8]), .C(n2209), .Y(\U3/U9/Z_8 ) );
  and2a3 U2480 ( .A(n2208), .B(reg2[8]), .Y(n2209) );
  ao1a1 U2481 ( .A(n2206), .B(reg1[7]), .C(n2210), .Y(\U3/U9/Z_7 ) );
  and2a3 U2482 ( .A(n2208), .B(reg2[7]), .Y(n2210) );
  ao1a1 U2483 ( .A(n2206), .B(reg1[6]), .C(n2211), .Y(\U3/U9/Z_6 ) );
  and2a3 U2484 ( .A(n2208), .B(reg2[6]), .Y(n2211) );
  ao1a1 U2485 ( .A(n2206), .B(reg1[5]), .C(n2212), .Y(\U3/U9/Z_5 ) );
  and2a3 U2486 ( .A(n2208), .B(reg2[5]), .Y(n2212) );
  ao1a1 U2487 ( .A(n2206), .B(reg1[4]), .C(n2213), .Y(\U3/U9/Z_4 ) );
  and2a3 U2488 ( .A(n2208), .B(reg2[4]), .Y(n2213) );
  or2a1 U2489 ( .A(\U3/U9/Z_31 ), .B(\U3/U10/Z_0 ), .Y(\U3/U9/Z_30 ) );
  ao1a1 U2490 ( .A(n2206), .B(reg1[19]), .C(n2214), .Y(\U3/U9/Z_31 ) );
  and2a3 U2491 ( .A(n2208), .B(reg2[19]), .Y(n2214) );
  ao1a1 U2492 ( .A(n2206), .B(reg1[3]), .C(n2215), .Y(\U3/U9/Z_3 ) );
  and2a3 U2493 ( .A(n2208), .B(reg2[3]), .Y(n2215) );
  ao1a1 U2494 ( .A(n2206), .B(reg1[2]), .C(n2216), .Y(\U3/U9/Z_2 ) );
  and2a3 U2495 ( .A(n2208), .B(reg2[2]), .Y(n2216) );
  ao1a1 U2496 ( .A(n2206), .B(reg1[18]), .C(n2217), .Y(\U3/U9/Z_18 ) );
  and2a3 U2497 ( .A(n2208), .B(reg2[18]), .Y(n2217) );
  ao1a1 U2498 ( .A(n2206), .B(reg1[17]), .C(n2218), .Y(\U3/U9/Z_17 ) );
  and2a3 U2499 ( .A(n2208), .B(reg2[17]), .Y(n2218) );
  ao1a1 U2500 ( .A(n2206), .B(reg1[16]), .C(n2219), .Y(\U3/U9/Z_16 ) );
  and2a3 U2501 ( .A(n2208), .B(reg2[16]), .Y(n2219) );
  ao1a1 U2502 ( .A(n2206), .B(reg1[15]), .C(n2220), .Y(\U3/U9/Z_15 ) );
  and2a3 U2503 ( .A(n2208), .B(reg2[15]), .Y(n2220) );
  ao1a1 U2504 ( .A(n2206), .B(reg1[14]), .C(n2221), .Y(\U3/U9/Z_14 ) );
  and2a3 U2505 ( .A(n2208), .B(reg2[14]), .Y(n2221) );
  ao1a1 U2506 ( .A(n2206), .B(reg1[13]), .C(n2222), .Y(\U3/U9/Z_13 ) );
  and2a3 U2507 ( .A(n2208), .B(reg2[13]), .Y(n2222) );
  ao1a1 U2508 ( .A(n2206), .B(reg1[12]), .C(n2223), .Y(\U3/U9/Z_12 ) );
  and2a3 U2509 ( .A(n2208), .B(reg2[12]), .Y(n2223) );
  ao1a1 U2510 ( .A(n2206), .B(reg1[11]), .C(n2224), .Y(\U3/U9/Z_11 ) );
  and2a3 U2511 ( .A(n2208), .B(reg2[11]), .Y(n2224) );
  ao1a1 U2512 ( .A(n2206), .B(reg1[10]), .C(n2225), .Y(\U3/U9/Z_10 ) );
  and2a3 U2513 ( .A(n2208), .B(reg2[10]), .Y(n2225) );
  ao1a1 U2514 ( .A(n2206), .B(reg1[1]), .C(n2226), .Y(\U3/U9/Z_1 ) );
  and2a3 U2515 ( .A(n2208), .B(reg2[1]), .Y(n2226) );
  or3a1 U2516 ( .A(n2227), .B(n2228), .C(n2229), .Y(\U3/U9/Z_0 ) );
  and2a3 U2517 ( .A(reg1[0]), .B(n2206), .Y(n2229) );
  and2a3 U2518 ( .A(reg2[0]), .B(n2208), .Y(n2228) );
  and3a1 U2519 ( .A(N654), .B(N685), .C(n2230), .Y(n2227) );
  or3a1 U2520 ( .A(n2231), .B(n2232), .C(n2233), .Y(\U3/U8/Z_9 ) );
  and2a3 U2521 ( .A(\U3/U10/Z_0 ), .B(N663), .Y(n2233) );
  and2a3 U2522 ( .A(n2230), .B(N664), .Y(n2231) );
  or3a1 U2523 ( .A(n2235), .B(n2236), .C(n2237), .Y(\U3/U8/Z_8 ) );
  and2a3 U2524 ( .A(\U3/U10/Z_0 ), .B(N662), .Y(n2237) );
  and2a3 U2525 ( .A(n2230), .B(N663), .Y(n2235) );
  or3a1 U2526 ( .A(n2238), .B(n2239), .C(n2240), .Y(\U3/U8/Z_7 ) );
  and2a3 U2527 ( .A(\U3/U10/Z_0 ), .B(N661), .Y(n2240) );
  and2a3 U2528 ( .A(n2230), .B(N662), .Y(n2238) );
  or3a1 U2529 ( .A(n2241), .B(n2242), .C(n2243), .Y(\U3/U8/Z_6 ) );
  and2a3 U2530 ( .A(\U3/U10/Z_0 ), .B(N660), .Y(n2243) );
  and2a3 U2531 ( .A(N549), .B(n2234), .Y(n2242) );
  and2a3 U2532 ( .A(n2230), .B(N661), .Y(n2241) );
  or3a1 U2533 ( .A(n2244), .B(n2245), .C(n2246), .Y(\U3/U8/Z_5 ) );
  and2a3 U2534 ( .A(\U3/U10/Z_0 ), .B(N659), .Y(n2246) );
  and2a3 U2535 ( .A(n2230), .B(N660), .Y(n2244) );
  or3a1 U2536 ( .A(n2247), .B(n2248), .C(n2249), .Y(\U3/U8/Z_4 ) );
  and2a3 U2537 ( .A(\U3/U10/Z_0 ), .B(N658), .Y(n2249) );
  and2a3 U2538 ( .A(n2230), .B(N659), .Y(n2247) );
  or2a1 U2539 ( .A(\U3/U10/Z_0 ), .B(\U3/U8/Z_31 ), .Y(\U3/U8/Z_30 ) );
  ao1a1 U2540 ( .A(N685), .B(n2230), .C(n2250), .Y(\U3/U8/Z_31 ) );
  or3a1 U2541 ( .A(n2251), .B(n2252), .C(n2253), .Y(\U3/U8/Z_3 ) );
  and2a3 U2542 ( .A(\U3/U10/Z_0 ), .B(N657), .Y(n2253) );
  and2a3 U2543 ( .A(n2230), .B(N658), .Y(n2251) );
  ao1f1 U2544 ( .A(n2254), .B(n2255), .C(n2256), .Y(\U3/U8/Z_29 ) );
  oa1f1 U2545 ( .A(n2230), .B(N684), .C(n2250), .Y(n2256) );
  ao1f1 U2546 ( .A(n2257), .B(n2255), .C(n2258), .Y(\U3/U8/Z_28 ) );
  oa1f1 U2547 ( .A(n2230), .B(N683), .C(n2250), .Y(n2258) );
  ao1f1 U2548 ( .A(n2259), .B(n2255), .C(n2260), .Y(\U3/U8/Z_27 ) );
  oa1f1 U2549 ( .A(n2230), .B(N682), .C(n2250), .Y(n2260) );
  ao1f1 U2550 ( .A(n2261), .B(n2255), .C(n2262), .Y(\U3/U8/Z_26 ) );
  oa1f1 U2551 ( .A(n2230), .B(N681), .C(n2250), .Y(n2262) );
  ao1f1 U2552 ( .A(n2263), .B(n2255), .C(n2264), .Y(\U3/U8/Z_25 ) );
  oa1f1 U2553 ( .A(n2230), .B(N680), .C(n2250), .Y(n2264) );
  ao1f1 U2554 ( .A(n2265), .B(n2255), .C(n2266), .Y(\U3/U8/Z_24 ) );
  oa1f1 U2555 ( .A(n2230), .B(N679), .C(n2250), .Y(n2266) );
  ao1f1 U2556 ( .A(n2267), .B(n2255), .C(n2268), .Y(\U3/U8/Z_23 ) );
  oa1f1 U2557 ( .A(n2230), .B(N678), .C(n2250), .Y(n2268) );
  ao1f1 U2558 ( .A(n2269), .B(n2255), .C(n2270), .Y(\U3/U8/Z_22 ) );
  oa1f1 U2559 ( .A(n2230), .B(N677), .C(n2250), .Y(n2270) );
  ao1f1 U2560 ( .A(n2271), .B(n2255), .C(n2272), .Y(\U3/U8/Z_21 ) );
  oa1f1 U2561 ( .A(n2230), .B(N676), .C(n2250), .Y(n2272) );
  ao1f1 U2562 ( .A(n2273), .B(n2255), .C(n2274), .Y(\U3/U8/Z_20 ) );
  oa1f1 U2563 ( .A(n2230), .B(N675), .C(n2250), .Y(n2274) );
  or3a1 U2564 ( .A(n2275), .B(n2276), .C(n2277), .Y(\U3/U8/Z_2 ) );
  and2a3 U2565 ( .A(\U3/U10/Z_0 ), .B(N656), .Y(n2277) );
  and2a3 U2566 ( .A(N553), .B(n2234), .Y(n2276) );
  and2a3 U2567 ( .A(n2230), .B(N657), .Y(n2275) );
  ao1f1 U2568 ( .A(n2278), .B(n2255), .C(n2279), .Y(\U3/U8/Z_19 ) );
  oa1f1 U2569 ( .A(n2230), .B(N674), .C(n2250), .Y(n2279) );
  and2a3 U2570 ( .A(n2234), .B(N536), .Y(n2250) );
  or3a1 U2571 ( .A(n2280), .B(n2281), .C(n2282), .Y(\U3/U8/Z_18 ) );
  and2a3 U2572 ( .A(\U3/U10/Z_0 ), .B(N672), .Y(n2282) );
  and2a3 U2573 ( .A(N537), .B(n2234), .Y(n2281) );
  and2a3 U2574 ( .A(n2230), .B(N673), .Y(n2280) );
  or3a1 U2575 ( .A(n2283), .B(n2284), .C(n2285), .Y(\U3/U8/Z_17 ) );
  and2a3 U2576 ( .A(\U3/U10/Z_0 ), .B(N671), .Y(n2285) );
  and2a3 U2577 ( .A(N538), .B(n2234), .Y(n2284) );
  and2a3 U2578 ( .A(n2230), .B(N672), .Y(n2283) );
  or3a1 U2579 ( .A(n2286), .B(n2287), .C(n2288), .Y(\U3/U8/Z_16 ) );
  and2a3 U2580 ( .A(\U3/U10/Z_0 ), .B(N670), .Y(n2288) );
  and2a3 U2581 ( .A(N539), .B(n2234), .Y(n2287) );
  and2a3 U2582 ( .A(n2230), .B(N671), .Y(n2286) );
  or3a1 U2583 ( .A(n2289), .B(n2290), .C(n2291), .Y(\U3/U8/Z_15 ) );
  and2a3 U2584 ( .A(\U3/U10/Z_0 ), .B(N669), .Y(n2291) );
  and2a3 U2585 ( .A(N540), .B(n2234), .Y(n2290) );
  and2a3 U2586 ( .A(n2230), .B(N670), .Y(n2289) );
  or3a1 U2587 ( .A(n2292), .B(n2293), .C(n2294), .Y(\U3/U8/Z_14 ) );
  and2a3 U2588 ( .A(\U3/U10/Z_0 ), .B(N668), .Y(n2294) );
  and2a3 U2589 ( .A(N541), .B(n2234), .Y(n2293) );
  and2a3 U2590 ( .A(n2230), .B(N669), .Y(n2292) );
  or3a1 U2591 ( .A(n2295), .B(n2296), .C(n2297), .Y(\U3/U8/Z_13 ) );
  and2a3 U2592 ( .A(\U3/U10/Z_0 ), .B(N667), .Y(n2297) );
  and2a3 U2593 ( .A(N542), .B(n2234), .Y(n2296) );
  and2a3 U2594 ( .A(n2230), .B(N668), .Y(n2295) );
  or3a1 U2595 ( .A(n2298), .B(n2299), .C(n2300), .Y(\U3/U8/Z_12 ) );
  and2a3 U2596 ( .A(\U3/U10/Z_0 ), .B(N666), .Y(n2300) );
  and2a3 U2597 ( .A(N543), .B(n2234), .Y(n2299) );
  and2a3 U2598 ( .A(n2230), .B(N667), .Y(n2298) );
  or3a1 U2599 ( .A(n2301), .B(n2302), .C(n2303), .Y(\U3/U8/Z_11 ) );
  and2a3 U2600 ( .A(\U3/U10/Z_0 ), .B(N665), .Y(n2303) );
  and2a3 U2601 ( .A(N544), .B(n2234), .Y(n2302) );
  and2a3 U2602 ( .A(n2230), .B(N666), .Y(n2301) );
  or3a1 U2603 ( .A(n2304), .B(n2305), .C(n2306), .Y(\U3/U8/Z_10 ) );
  and2a3 U2604 ( .A(\U3/U10/Z_0 ), .B(N664), .Y(n2306) );
  and2a3 U2605 ( .A(N545), .B(n2234), .Y(n2305) );
  and2a3 U2606 ( .A(n2230), .B(N665), .Y(n2304) );
  or3a1 U2607 ( .A(n2307), .B(n2308), .C(n2309), .Y(\U3/U8/Z_1 ) );
  and2a3 U2608 ( .A(\U3/U10/Z_0 ), .B(N655), .Y(n2309) );
  and2a3 U2609 ( .A(N554), .B(n2234), .Y(n2308) );
  and2a3 U2610 ( .A(n2230), .B(N656), .Y(n2307) );
  or3a1 U2611 ( .A(n2310), .B(n2311), .C(n2312), .Y(\U3/U8/Z_0 ) );
  and2a3 U2612 ( .A(\U3/U10/Z_0 ), .B(N654), .Y(n2312) );
  and2a3 U2613 ( .A(N555), .B(n2234), .Y(n2311) );
  and2a3 U2614 ( .A(n2230), .B(N655), .Y(n2310) );
  ao1f1 U2615 ( .A(n2318), .B(n2319), .C(n2320), .Y(\U3/U7/Z_9 ) );
  or2a1 U2616 ( .A(n2321), .B(n2322), .Y(n2320) );
  ao1f1 U2617 ( .A(n2323), .B(n2319), .C(n2324), .Y(\U3/U7/Z_8 ) );
  or2a1 U2618 ( .A(n2325), .B(n2322), .Y(n2324) );
  ao1f1 U2619 ( .A(n2326), .B(n2319), .C(n2327), .Y(\U3/U7/Z_7 ) );
  or2a1 U2620 ( .A(n2328), .B(n2322), .Y(n2327) );
  ao1f1 U2621 ( .A(n2329), .B(n2319), .C(n2330), .Y(\U3/U7/Z_6 ) );
  or2a1 U2622 ( .A(n2331), .B(n2322), .Y(n2330) );
  ao1f1 U2623 ( .A(n2332), .B(n2319), .C(n2333), .Y(\U3/U7/Z_5 ) );
  or2a1 U2624 ( .A(n2334), .B(n2322), .Y(n2333) );
  ao1f1 U2625 ( .A(n2335), .B(n2319), .C(n2336), .Y(\U3/U7/Z_4 ) );
  or2a1 U2626 ( .A(n2337), .B(n2322), .Y(n2336) );
  and2a3 U2627 ( .A(N970), .B(n2338), .Y(\U3/U7/Z_31 ) );
  and2a3 U2628 ( .A(N969), .B(n2338), .Y(\U3/U7/Z_30 ) );
  ao1f1 U2629 ( .A(n2339), .B(n2319), .C(n2340), .Y(\U3/U7/Z_3 ) );
  or2a1 U2630 ( .A(n2341), .B(n2322), .Y(n2340) );
  ao1f1 U2631 ( .A(n2319), .B(n2342), .C(n2343), .Y(\U3/U7/Z_29 ) );
  or2a1 U2632 ( .A(n2257), .B(n2322), .Y(n2343) );
  ao1f1 U2633 ( .A(n2319), .B(n2344), .C(n2345), .Y(\U3/U7/Z_28 ) );
  or2a1 U2634 ( .A(n2259), .B(n2322), .Y(n2345) );
  ao1f1 U2635 ( .A(n2319), .B(n2346), .C(n2347), .Y(\U3/U7/Z_27 ) );
  or2a1 U2636 ( .A(n2261), .B(n2322), .Y(n2347) );
  ao1f1 U2637 ( .A(n2319), .B(n2348), .C(n2349), .Y(\U3/U7/Z_26 ) );
  or2a1 U2638 ( .A(n2263), .B(n2322), .Y(n2349) );
  ao1f1 U2639 ( .A(n2319), .B(n2350), .C(n2351), .Y(\U3/U7/Z_25 ) );
  or2a1 U2640 ( .A(n2265), .B(n2322), .Y(n2351) );
  ao1f1 U2641 ( .A(n2319), .B(n2352), .C(n2353), .Y(\U3/U7/Z_24 ) );
  or2a1 U2642 ( .A(n2267), .B(n2322), .Y(n2353) );
  ao1f1 U2643 ( .A(n2319), .B(n2354), .C(n2355), .Y(\U3/U7/Z_23 ) );
  or2a1 U2644 ( .A(n2269), .B(n2322), .Y(n2355) );
  ao1f1 U2645 ( .A(n2319), .B(n2356), .C(n2357), .Y(\U3/U7/Z_22 ) );
  or2a1 U2646 ( .A(n2271), .B(n2322), .Y(n2357) );
  ao1f1 U2647 ( .A(n2319), .B(n2358), .C(n2359), .Y(\U3/U7/Z_21 ) );
  or2a1 U2648 ( .A(n2273), .B(n2322), .Y(n2359) );
  ao1f1 U2649 ( .A(n2319), .B(n2360), .C(n2361), .Y(\U3/U7/Z_20 ) );
  or2a1 U2650 ( .A(n2278), .B(n2322), .Y(n2361) );
  ao1f1 U2651 ( .A(n2362), .B(n2319), .C(n2363), .Y(\U3/U7/Z_2 ) );
  or2a1 U2652 ( .A(n2364), .B(n2322), .Y(n2363) );
  ao1f1 U2653 ( .A(n2365), .B(n2319), .C(n2366), .Y(\U3/U7/Z_19 ) );
  or2a1 U2654 ( .A(n2367), .B(n2322), .Y(n2366) );
  ao1f1 U2655 ( .A(n2368), .B(n2319), .C(n2369), .Y(\U3/U7/Z_18 ) );
  or2a1 U2656 ( .A(n2370), .B(n2322), .Y(n2369) );
  ao1f1 U2657 ( .A(n2371), .B(n2319), .C(n2372), .Y(\U3/U7/Z_17 ) );
  or2a1 U2658 ( .A(n2373), .B(n2322), .Y(n2372) );
  ao1f1 U2659 ( .A(n2374), .B(n2319), .C(n2375), .Y(\U3/U7/Z_16 ) );
  or2a1 U2660 ( .A(n2376), .B(n2322), .Y(n2375) );
  ao1f1 U2661 ( .A(n2377), .B(n2319), .C(n2378), .Y(\U3/U7/Z_15 ) );
  or2a1 U2662 ( .A(n2379), .B(n2322), .Y(n2378) );
  ao1f1 U2663 ( .A(n2380), .B(n2319), .C(n2381), .Y(\U3/U7/Z_14 ) );
  or2a1 U2664 ( .A(n2382), .B(n2322), .Y(n2381) );
  ao1f1 U2665 ( .A(n2383), .B(n2319), .C(n2384), .Y(\U3/U7/Z_13 ) );
  or2a1 U2666 ( .A(n2385), .B(n2322), .Y(n2384) );
  ao1f1 U2667 ( .A(n2386), .B(n2319), .C(n2387), .Y(\U3/U7/Z_12 ) );
  or2a1 U2668 ( .A(n2388), .B(n2322), .Y(n2387) );
  ao1f1 U2669 ( .A(n2389), .B(n2319), .C(n2390), .Y(\U3/U7/Z_11 ) );
  or2a1 U2670 ( .A(n2391), .B(n2322), .Y(n2390) );
  ao1f1 U2671 ( .A(n2392), .B(n2319), .C(n2393), .Y(\U3/U7/Z_10 ) );
  or2a1 U2672 ( .A(n2394), .B(n2322), .Y(n2393) );
  ao1f1 U2673 ( .A(n2395), .B(n2319), .C(n2396), .Y(\U3/U7/Z_1 ) );
  or2a1 U2674 ( .A(n2397), .B(n2322), .Y(n2396) );
  and2a3 U2675 ( .A(n2338), .B(N939), .Y(\U3/U7/Z_0 ) );
  ao1f1 U2676 ( .A(n2255), .B(n2398), .C(n2399), .Y(\U3/U6/Z_9 ) );
  oa1f1 U2677 ( .A(n2400), .B(N663), .C(n2401), .Y(n2399) );
  ao1f1 U2678 ( .A(n2255), .B(n2402), .C(n2403), .Y(\U3/U6/Z_8 ) );
  oa1f1 U2679 ( .A(n2400), .B(N662), .C(n2401), .Y(n2403) );
  ao1f1 U2680 ( .A(n2255), .B(n2404), .C(n2405), .Y(\U3/U6/Z_7 ) );
  oa1f1 U2681 ( .A(n2400), .B(N661), .C(n2401), .Y(n2405) );
  ao1f1 U2682 ( .A(n2255), .B(n2406), .C(n2407), .Y(\U3/U6/Z_6 ) );
  oa1f1 U2683 ( .A(n2400), .B(N660), .C(n2401), .Y(n2407) );
  ao1f1 U2684 ( .A(n2255), .B(n2408), .C(n2409), .Y(\U3/U6/Z_5 ) );
  oa1f1 U2685 ( .A(n2400), .B(N659), .C(n2401), .Y(n2409) );
  ao1f1 U2686 ( .A(n2255), .B(n2410), .C(n2411), .Y(\U3/U6/Z_4 ) );
  oa1f1 U2687 ( .A(n2400), .B(N658), .C(n2401), .Y(n2411) );
  ao1a1 U2688 ( .A(N685), .B(n2400), .C(n2412), .Y(\U3/U6/Z_31 ) );
  and2a3 U2689 ( .A(\U3/U10/Z_0 ), .B(n189), .Y(n2412) );
  ao1a1 U2690 ( .A(N684), .B(n2400), .C(n2413), .Y(\U3/U6/Z_30 ) );
  and2a3 U2691 ( .A(\U3/U10/Z_0 ), .B(n190), .Y(n2413) );
  ao1f1 U2692 ( .A(n2255), .B(n2414), .C(n2415), .Y(\U3/U6/Z_3 ) );
  oa1f1 U2693 ( .A(n2400), .B(N657), .C(n2401), .Y(n2415) );
  ao1f1 U2694 ( .A(n2255), .B(n2416), .C(n2417), .Y(\U3/U6/Z_29 ) );
  oa1f1 U2695 ( .A(n2400), .B(N683), .C(n2401), .Y(n2417) );
  ao1f1 U2696 ( .A(n2255), .B(n2418), .C(n2419), .Y(\U3/U6/Z_28 ) );
  oa1f1 U2697 ( .A(n2400), .B(N682), .C(n2401), .Y(n2419) );
  ao1f1 U2698 ( .A(n2255), .B(n2420), .C(n2421), .Y(\U3/U6/Z_27 ) );
  oa1f1 U2699 ( .A(n2400), .B(N681), .C(n2401), .Y(n2421) );
  ao1f1 U2700 ( .A(n2255), .B(n2422), .C(n2423), .Y(\U3/U6/Z_26 ) );
  oa1f1 U2701 ( .A(n2400), .B(N680), .C(n2401), .Y(n2423) );
  ao1f1 U2702 ( .A(n2255), .B(n2424), .C(n2425), .Y(\U3/U6/Z_25 ) );
  oa1f1 U2703 ( .A(n2400), .B(N679), .C(n2401), .Y(n2425) );
  ao1f1 U2704 ( .A(n2255), .B(n2426), .C(n2427), .Y(\U3/U6/Z_24 ) );
  oa1f1 U2705 ( .A(n2400), .B(N678), .C(n2401), .Y(n2427) );
  ao1f1 U2706 ( .A(n2255), .B(n2428), .C(n2429), .Y(\U3/U6/Z_23 ) );
  oa1f1 U2707 ( .A(n2400), .B(N677), .C(n2401), .Y(n2429) );
  ao1f1 U2708 ( .A(n2255), .B(n2430), .C(n2431), .Y(\U3/U6/Z_22 ) );
  oa1f1 U2709 ( .A(n2400), .B(N676), .C(n2401), .Y(n2431) );
  ao1f1 U2710 ( .A(n2255), .B(n2432), .C(n2433), .Y(\U3/U6/Z_21 ) );
  oa1f1 U2711 ( .A(n2400), .B(N675), .C(n2401), .Y(n2433) );
  ao1f1 U2712 ( .A(n2255), .B(n2434), .C(n2435), .Y(\U3/U6/Z_20 ) );
  oa1f1 U2713 ( .A(n2400), .B(N674), .C(n2401), .Y(n2435) );
  ao1f1 U2714 ( .A(n2255), .B(n2436), .C(n2437), .Y(\U3/U6/Z_2 ) );
  oa1f1 U2715 ( .A(n2400), .B(N656), .C(n2401), .Y(n2437) );
  ao1f1 U2716 ( .A(n2255), .B(n2438), .C(n2439), .Y(\U3/U6/Z_19 ) );
  oa1f1 U2717 ( .A(n2400), .B(N673), .C(n2401), .Y(n2439) );
  ao1f1 U2718 ( .A(n2255), .B(n2440), .C(n2441), .Y(\U3/U6/Z_18 ) );
  oa1f1 U2719 ( .A(n2400), .B(N672), .C(n2401), .Y(n2441) );
  ao1f1 U2720 ( .A(n2255), .B(n2442), .C(n2443), .Y(\U3/U6/Z_17 ) );
  oa1f1 U2721 ( .A(n2400), .B(N671), .C(n2401), .Y(n2443) );
  ao1f1 U2722 ( .A(n2255), .B(n2444), .C(n2445), .Y(\U3/U6/Z_16 ) );
  oa1f1 U2723 ( .A(n2400), .B(N670), .C(n2401), .Y(n2445) );
  ao1f1 U2724 ( .A(n2255), .B(n2446), .C(n2447), .Y(\U3/U6/Z_15 ) );
  oa1f1 U2725 ( .A(n2400), .B(N669), .C(n2401), .Y(n2447) );
  ao1f1 U2726 ( .A(n2255), .B(n2448), .C(n2449), .Y(\U3/U6/Z_14 ) );
  oa1f1 U2727 ( .A(n2400), .B(N668), .C(n2401), .Y(n2449) );
  ao1f1 U2728 ( .A(n2255), .B(n2450), .C(n2451), .Y(\U3/U6/Z_13 ) );
  oa1f1 U2729 ( .A(n2400), .B(N667), .C(n2401), .Y(n2451) );
  ao1f1 U2730 ( .A(n2255), .B(n2452), .C(n2453), .Y(\U3/U6/Z_12 ) );
  oa1f1 U2731 ( .A(n2400), .B(N666), .C(n2401), .Y(n2453) );
  ao1f1 U2732 ( .A(n2255), .B(n2454), .C(n2455), .Y(\U3/U6/Z_11 ) );
  oa1f1 U2733 ( .A(n2400), .B(N665), .C(n2401), .Y(n2455) );
  ao1f1 U2734 ( .A(n2255), .B(n2456), .C(n2457), .Y(\U3/U6/Z_10 ) );
  oa1f1 U2735 ( .A(n2400), .B(N664), .C(n2401), .Y(n2457) );
  ao1f1 U2736 ( .A(n2255), .B(n2458), .C(n2459), .Y(\U3/U6/Z_1 ) );
  oa1f1 U2737 ( .A(n2400), .B(N655), .C(n2401), .Y(n2459) );
  ao1f1 U2738 ( .A(n2255), .B(n2460), .C(n2461), .Y(\U3/U6/Z_0 ) );
  oa1f1 U2739 ( .A(n2400), .B(N654), .C(n2401), .Y(n2461) );
  inv1a1 U2740 ( .A(n2466), .Y(n2465) );
  inv1a1 U2741 ( .A(n220), .Y(n2460) );
  or3a1 U2742 ( .A(n2467), .B(n2468), .C(n2469), .Y(\U3/U4/Z_9 ) );
  and2a3 U2743 ( .A(reg1[9]), .B(n2470), .Y(n2469) );
  and2a3 U2744 ( .A(reg2[9]), .B(n2471), .Y(n2468) );
  and2a3 U2745 ( .A(n2472), .B(N948), .Y(n2467) );
  or3a1 U2746 ( .A(n2473), .B(n2474), .C(n2475), .Y(\U3/U4/Z_8 ) );
  and2a3 U2747 ( .A(reg1[8]), .B(n2470), .Y(n2475) );
  and2a3 U2748 ( .A(reg2[8]), .B(n2471), .Y(n2474) );
  and2a3 U2749 ( .A(n2472), .B(N947), .Y(n2473) );
  or3a1 U2750 ( .A(n2476), .B(n2477), .C(n2478), .Y(\U3/U4/Z_7 ) );
  and2a3 U2751 ( .A(reg1[7]), .B(n2470), .Y(n2478) );
  and2a3 U2752 ( .A(reg2[7]), .B(n2471), .Y(n2477) );
  and2a3 U2753 ( .A(n2472), .B(N946), .Y(n2476) );
  or3a1 U2754 ( .A(n2479), .B(n2480), .C(n2481), .Y(\U3/U4/Z_6 ) );
  and2a3 U2755 ( .A(reg1[6]), .B(n2470), .Y(n2481) );
  and2a3 U2756 ( .A(reg2[6]), .B(n2471), .Y(n2480) );
  and2a3 U2757 ( .A(n2472), .B(N945), .Y(n2479) );
  or3a1 U2758 ( .A(n2482), .B(n2483), .C(n2484), .Y(\U3/U4/Z_5 ) );
  and2a3 U2759 ( .A(reg1[5]), .B(n2470), .Y(n2484) );
  and2a3 U2760 ( .A(reg2[5]), .B(n2471), .Y(n2483) );
  and2a3 U2761 ( .A(n2472), .B(N944), .Y(n2482) );
  or3a1 U2762 ( .A(n2485), .B(n2486), .C(n2487), .Y(\U3/U4/Z_4 ) );
  and2a3 U2763 ( .A(reg1[4]), .B(n2470), .Y(n2487) );
  and2a3 U2764 ( .A(reg2[4]), .B(n2471), .Y(n2486) );
  and2a3 U2765 ( .A(n2472), .B(N943), .Y(n2485) );
  or3a1 U2766 ( .A(n2488), .B(n2489), .C(n2490), .Y(\U3/U4/Z_3 ) );
  and2a3 U2767 ( .A(reg1[3]), .B(n2470), .Y(n2490) );
  and2a3 U2768 ( .A(reg2[3]), .B(n2471), .Y(n2489) );
  and2a3 U2769 ( .A(n2472), .B(N942), .Y(n2488) );
  ao1f1 U2770 ( .A(n2491), .B(n2344), .C(n2492), .Y(\U3/U4/Z_28 ) );
  ao1f1 U2771 ( .A(n2491), .B(n2346), .C(n2492), .Y(\U3/U4/Z_27 ) );
  ao1f1 U2772 ( .A(n2491), .B(n2348), .C(n2492), .Y(\U3/U4/Z_26 ) );
  ao1f1 U2773 ( .A(n2491), .B(n2350), .C(n2492), .Y(\U3/U4/Z_25 ) );
  ao1f1 U2774 ( .A(n2491), .B(n2352), .C(n2492), .Y(\U3/U4/Z_24 ) );
  ao1f1 U2775 ( .A(n2491), .B(n2354), .C(n2492), .Y(\U3/U4/Z_23 ) );
  ao1f1 U2776 ( .A(n2491), .B(n2356), .C(n2492), .Y(\U3/U4/Z_22 ) );
  ao1f1 U2777 ( .A(n2491), .B(n2358), .C(n2492), .Y(\U3/U4/Z_21 ) );
  ao1f1 U2778 ( .A(n2491), .B(n2360), .C(n2492), .Y(\U3/U4/Z_20 ) );
  or3a1 U2779 ( .A(n2493), .B(n2494), .C(n2495), .Y(\U3/U4/Z_2 ) );
  and2a3 U2780 ( .A(reg1[2]), .B(n2470), .Y(n2495) );
  and2a3 U2781 ( .A(reg2[2]), .B(n2471), .Y(n2494) );
  and2a3 U2782 ( .A(n2472), .B(N941), .Y(n2493) );
  ao1f1 U2783 ( .A(n2365), .B(n2491), .C(n2492), .Y(\U3/U4/Z_19 ) );
  and2a3 U2784 ( .A(n2470), .B(reg1[19]), .Y(n2496) );
  or3a1 U2785 ( .A(n2497), .B(n2498), .C(n2499), .Y(\U3/U4/Z_18 ) );
  and2a3 U2786 ( .A(reg1[18]), .B(n2470), .Y(n2499) );
  and2a3 U2787 ( .A(reg2[18]), .B(n2471), .Y(n2498) );
  and2a3 U2788 ( .A(n2472), .B(N957), .Y(n2497) );
  or3a1 U2789 ( .A(n2500), .B(n2501), .C(n2502), .Y(\U3/U4/Z_17 ) );
  and2a3 U2790 ( .A(reg1[17]), .B(n2470), .Y(n2502) );
  and2a3 U2791 ( .A(reg2[17]), .B(n2471), .Y(n2501) );
  and2a3 U2792 ( .A(n2472), .B(N956), .Y(n2500) );
  or3a1 U2793 ( .A(n2503), .B(n2504), .C(n2505), .Y(\U3/U4/Z_16 ) );
  and2a3 U2794 ( .A(reg1[16]), .B(n2470), .Y(n2505) );
  and2a3 U2795 ( .A(reg2[16]), .B(n2471), .Y(n2504) );
  and2a3 U2796 ( .A(n2472), .B(N955), .Y(n2503) );
  or3a1 U2797 ( .A(n2506), .B(n2507), .C(n2508), .Y(\U3/U4/Z_15 ) );
  and2a3 U2798 ( .A(reg1[15]), .B(n2470), .Y(n2508) );
  and2a3 U2799 ( .A(reg2[15]), .B(n2471), .Y(n2507) );
  and2a3 U2800 ( .A(n2472), .B(N954), .Y(n2506) );
  or3a1 U2801 ( .A(n2509), .B(n2510), .C(n2511), .Y(\U3/U4/Z_14 ) );
  and2a3 U2802 ( .A(reg1[14]), .B(n2470), .Y(n2511) );
  and2a3 U2803 ( .A(reg2[14]), .B(n2471), .Y(n2510) );
  and2a3 U2804 ( .A(n2472), .B(N953), .Y(n2509) );
  or3a1 U2805 ( .A(n2512), .B(n2513), .C(n2514), .Y(\U3/U4/Z_13 ) );
  and2a3 U2806 ( .A(reg1[13]), .B(n2470), .Y(n2514) );
  and2a3 U2807 ( .A(reg2[13]), .B(n2471), .Y(n2513) );
  and2a3 U2808 ( .A(n2472), .B(N952), .Y(n2512) );
  or3a1 U2809 ( .A(n2515), .B(n2516), .C(n2517), .Y(\U3/U4/Z_12 ) );
  and2a3 U2810 ( .A(reg1[12]), .B(n2470), .Y(n2517) );
  and2a3 U2811 ( .A(reg2[12]), .B(n2471), .Y(n2516) );
  and2a3 U2812 ( .A(n2472), .B(N951), .Y(n2515) );
  or3a1 U2813 ( .A(n2518), .B(n2519), .C(n2520), .Y(\U3/U4/Z_11 ) );
  and2a3 U2814 ( .A(reg1[11]), .B(n2470), .Y(n2520) );
  and2a3 U2815 ( .A(reg2[11]), .B(n2471), .Y(n2519) );
  and2a3 U2816 ( .A(n2472), .B(N950), .Y(n2518) );
  or3a1 U2817 ( .A(n2521), .B(n2522), .C(n2523), .Y(\U3/U4/Z_10 ) );
  and2a3 U2818 ( .A(reg1[10]), .B(n2470), .Y(n2523) );
  and2a3 U2819 ( .A(reg2[10]), .B(n2471), .Y(n2522) );
  and2a3 U2820 ( .A(n2472), .B(N949), .Y(n2521) );
  or3a1 U2821 ( .A(n2524), .B(n2525), .C(n2526), .Y(\U3/U4/Z_1 ) );
  and2a3 U2822 ( .A(reg1[1]), .B(n2470), .Y(n2526) );
  and2a3 U2823 ( .A(reg2[1]), .B(n2471), .Y(n2525) );
  and2a3 U2824 ( .A(n2472), .B(N940), .Y(n2524) );
  or3a1 U2825 ( .A(n2527), .B(n2528), .C(n2529), .Y(\U3/U4/Z_0 ) );
  and2a3 U2826 ( .A(reg1[0]), .B(n2470), .Y(n2529) );
  and2a3 U2827 ( .A(reg2[0]), .B(n2471), .Y(n2528) );
  and2a3 U2828 ( .A(n2472), .B(N939), .Y(n2527) );
  or2a1 U2829 ( .A(n2534), .B(n2535), .Y(n2533) );
  ao1f1 U2830 ( .A(n2536), .B(n2537), .C(n2538), .Y(\U3/U3/Z_9 ) );
  or2a1 U2831 ( .A(n2539), .B(n2394), .Y(n2538) );
  inv1a1 U2832 ( .A(N546), .Y(n2537) );
  ao1f1 U2833 ( .A(n2536), .B(n2540), .C(n2541), .Y(\U3/U3/Z_8 ) );
  or2a1 U2834 ( .A(n2539), .B(n2321), .Y(n2541) );
  inv1a1 U2835 ( .A(N547), .Y(n2540) );
  ao1f1 U2836 ( .A(n2536), .B(n2542), .C(n2543), .Y(\U3/U3/Z_7 ) );
  or2a1 U2837 ( .A(n2539), .B(n2325), .Y(n2543) );
  inv1a1 U2838 ( .A(N548), .Y(n2542) );
  ao1f1 U2839 ( .A(n2536), .B(n2544), .C(n2545), .Y(\U3/U3/Z_6 ) );
  or2a1 U2840 ( .A(n2539), .B(n2328), .Y(n2545) );
  inv1a1 U2841 ( .A(N549), .Y(n2544) );
  ao1f1 U2842 ( .A(n2536), .B(n2546), .C(n2547), .Y(\U3/U3/Z_5 ) );
  or2a1 U2843 ( .A(n2539), .B(n2331), .Y(n2547) );
  inv1a1 U2844 ( .A(N550), .Y(n2546) );
  ao1f1 U2845 ( .A(n2536), .B(n2548), .C(n2549), .Y(\U3/U3/Z_4 ) );
  or2a1 U2846 ( .A(n2539), .B(n2334), .Y(n2549) );
  inv1a1 U2847 ( .A(N551), .Y(n2548) );
  ao1f1 U2848 ( .A(n2536), .B(n2550), .C(n2551), .Y(\U3/U3/Z_3 ) );
  or2a1 U2849 ( .A(n2539), .B(n2337), .Y(n2551) );
  inv1a1 U2850 ( .A(N552), .Y(n2550) );
  ao1f1 U2851 ( .A(n2257), .B(n2539), .C(n2552), .Y(\U3/U3/Z_28 ) );
  ao1f1 U2852 ( .A(n2259), .B(n2539), .C(n2552), .Y(\U3/U3/Z_27 ) );
  ao1f1 U2853 ( .A(n2261), .B(n2539), .C(n2552), .Y(\U3/U3/Z_26 ) );
  ao1f1 U2854 ( .A(n2263), .B(n2539), .C(n2552), .Y(\U3/U3/Z_25 ) );
  ao1f1 U2855 ( .A(n2265), .B(n2539), .C(n2552), .Y(\U3/U3/Z_24 ) );
  ao1f1 U2856 ( .A(n2267), .B(n2539), .C(n2552), .Y(\U3/U3/Z_23 ) );
  ao1f1 U2857 ( .A(n2269), .B(n2539), .C(n2552), .Y(\U3/U3/Z_22 ) );
  ao1f1 U2858 ( .A(n2271), .B(n2539), .C(n2552), .Y(\U3/U3/Z_21 ) );
  ao1f1 U2859 ( .A(n2273), .B(n2539), .C(n2552), .Y(\U3/U3/Z_20 ) );
  ao1f1 U2860 ( .A(n2536), .B(n2553), .C(n2554), .Y(\U3/U3/Z_2 ) );
  or2a1 U2861 ( .A(n2539), .B(n2341), .Y(n2554) );
  inv1a1 U2862 ( .A(N553), .Y(n2553) );
  ao1f1 U2863 ( .A(n2539), .B(n2278), .C(n2552), .Y(\U3/U3/Z_19 ) );
  and2a3 U2864 ( .A(n2556), .B(N536), .Y(n2555) );
  ao1f1 U2865 ( .A(n2536), .B(n2557), .C(n2558), .Y(\U3/U3/Z_18 ) );
  or2a1 U2866 ( .A(n2539), .B(n2367), .Y(n2558) );
  inv1a1 U2867 ( .A(N537), .Y(n2557) );
  ao1f1 U2868 ( .A(n2536), .B(n2559), .C(n2560), .Y(\U3/U3/Z_17 ) );
  or2a1 U2869 ( .A(n2539), .B(n2370), .Y(n2560) );
  inv1a1 U2870 ( .A(N538), .Y(n2559) );
  ao1f1 U2871 ( .A(n2536), .B(n2561), .C(n2562), .Y(\U3/U3/Z_16 ) );
  or2a1 U2872 ( .A(n2539), .B(n2373), .Y(n2562) );
  inv1a1 U2873 ( .A(N539), .Y(n2561) );
  ao1f1 U2874 ( .A(n2536), .B(n2563), .C(n2564), .Y(\U3/U3/Z_15 ) );
  or2a1 U2875 ( .A(n2539), .B(n2376), .Y(n2564) );
  inv1a1 U2876 ( .A(N540), .Y(n2563) );
  ao1f1 U2877 ( .A(n2536), .B(n2565), .C(n2566), .Y(\U3/U3/Z_14 ) );
  or2a1 U2878 ( .A(n2539), .B(n2379), .Y(n2566) );
  inv1a1 U2879 ( .A(N541), .Y(n2565) );
  ao1f1 U2880 ( .A(n2536), .B(n2567), .C(n2568), .Y(\U3/U3/Z_13 ) );
  or2a1 U2881 ( .A(n2539), .B(n2382), .Y(n2568) );
  inv1a1 U2882 ( .A(N542), .Y(n2567) );
  ao1f1 U2883 ( .A(n2536), .B(n2569), .C(n2570), .Y(\U3/U3/Z_12 ) );
  or2a1 U2884 ( .A(n2539), .B(n2385), .Y(n2570) );
  inv1a1 U2885 ( .A(N543), .Y(n2569) );
  ao1f1 U2886 ( .A(n2536), .B(n2571), .C(n2572), .Y(\U3/U3/Z_11 ) );
  or2a1 U2887 ( .A(n2539), .B(n2388), .Y(n2572) );
  inv1a1 U2888 ( .A(N544), .Y(n2571) );
  ao1f1 U2889 ( .A(n2536), .B(n2573), .C(n2574), .Y(\U3/U3/Z_10 ) );
  or2a1 U2890 ( .A(n2539), .B(n2391), .Y(n2574) );
  inv1a1 U2891 ( .A(N545), .Y(n2573) );
  ao1f1 U2892 ( .A(n2536), .B(n2575), .C(n2576), .Y(\U3/U3/Z_1 ) );
  or2a1 U2893 ( .A(n2539), .B(n2364), .Y(n2576) );
  inv1a1 U2894 ( .A(N554), .Y(n2575) );
  ao1f1 U2895 ( .A(n2536), .B(n2577), .C(n2578), .Y(\U3/U3/Z_0 ) );
  or2a1 U2896 ( .A(n2539), .B(n2397), .Y(n2578) );
  or3a1 U2897 ( .A(n2535), .B(n2534), .C(n2530), .Y(n2579) );
  and2a3 U2898 ( .A(n2531), .B(n2580), .Y(n2530) );
  and2a3 U2899 ( .A(n2531), .B(n2581), .Y(n2534) );
  and2a3 U2900 ( .A(n2531), .B(n2582), .Y(n2535) );
  and2a3 U2901 ( .A(n2314), .B(n2583), .Y(n2531) );
  or2a1 U2902 ( .A(n2471), .B(n2470), .Y(n2556) );
  inv1a1 U2903 ( .A(n2588), .Y(n2585) );
  and2a3 U2904 ( .A(n2589), .B(n2314), .Y(n2588) );
  or2a1 U2905 ( .A(n2581), .B(n2593), .Y(n2591) );
  and2a3 U2906 ( .A(n2594), .B(N684), .Y(n2466) );
  inv1a1 U2907 ( .A(N685), .Y(n2594) );
  and2a3 U2908 ( .A(n2595), .B(N946), .Y(\U3/U1/Z_7 ) );
  and2a3 U2909 ( .A(n2595), .B(N942), .Y(\U3/U1/Z_3 ) );
  and2a3 U2910 ( .A(N967), .B(n2595), .Y(\U3/U1/Z_28 ) );
  and2a3 U2911 ( .A(N966), .B(n2595), .Y(\U3/U1/Z_27 ) );
  and2a3 U2912 ( .A(N965), .B(n2595), .Y(\U3/U1/Z_26 ) );
  and2a3 U2913 ( .A(N964), .B(n2595), .Y(\U3/U1/Z_25 ) );
  and2a3 U2914 ( .A(N963), .B(n2595), .Y(\U3/U1/Z_24 ) );
  and2a3 U2915 ( .A(N962), .B(n2595), .Y(\U3/U1/Z_23 ) );
  and2a3 U2916 ( .A(N961), .B(n2595), .Y(\U3/U1/Z_22 ) );
  and2a3 U2917 ( .A(N960), .B(n2595), .Y(\U3/U1/Z_21 ) );
  and2a3 U2918 ( .A(N959), .B(n2595), .Y(\U3/U1/Z_20 ) );
  and2a3 U2919 ( .A(n2595), .B(N954), .Y(\U3/U1/Z_15 ) );
  and2a3 U2920 ( .A(n2595), .B(N950), .Y(\U3/U1/Z_11 ) );
  and2a3 U2921 ( .A(n2595), .B(N940), .Y(\U3/U1/Z_1 ) );
  and2a3 U2922 ( .A(n2595), .B(N939), .Y(\U3/U1/Z_0 ) );
  and3a1 U2923 ( .A(n2599), .B(n2600), .C(n2601), .Y(n2598) );
  and2a3 U2924 ( .A(n2604), .B(n2596), .Y(n2601) );
  inv1a1 U2925 ( .A(n2600), .Y(n2603) );
  inv1a1 U2926 ( .A(n2602), .Y(n2599) );
  oa1f1 U2927 ( .A(n2605), .B(n2606), .C(N7058), .Y(N7124) );
  or3a1 U2928 ( .A(n2607), .B(n2463), .C(n2464), .Y(n2606) );
  and2a3 U2929 ( .A(n2596), .B(n2608), .Y(N7123) );
  mx2a1 U2930 ( .D0(datai[31]), .D1(N324), .S(state), .Y(N7057) );
  mx2a1 U2931 ( .D0(N323), .D1(datai[30]), .S(N7058), .Y(N7055) );
  mx2a1 U2932 ( .D0(N322), .D1(datai[29]), .S(N7058), .Y(N7053) );
  mx2a1 U2933 ( .D0(N321), .D1(datai[28]), .S(N7058), .Y(N7051) );
  mx2a1 U2934 ( .D0(N320), .D1(datai[27]), .S(N7058), .Y(N7049) );
  mx2a1 U2935 ( .D0(datai[26]), .D1(N319), .S(state), .Y(N7047) );
  mx2a1 U2936 ( .D0(datai[25]), .D1(N318), .S(state), .Y(N7045) );
  mx2a1 U2937 ( .D0(datai[24]), .D1(N317), .S(state), .Y(N7043) );
  mx2a1 U2938 ( .D0(datai[23]), .D1(N316), .S(state), .Y(N7041) );
  mx2a1 U2939 ( .D0(datai[22]), .D1(N315), .S(state), .Y(N7039) );
  mx2a1 U2940 ( .D0(datai[21]), .D1(N314), .S(state), .Y(N7037) );
  mx2a1 U2941 ( .D0(datai[20]), .D1(N313), .S(state), .Y(N7035) );
  mx2a1 U2942 ( .D0(datai[19]), .D1(N312), .S(state), .Y(N7033) );
  mx2a1 U2943 ( .D0(datai[18]), .D1(N311), .S(state), .Y(N7031) );
  mx2a1 U2944 ( .D0(datai[17]), .D1(N310), .S(state), .Y(N7029) );
  mx2a1 U2945 ( .D0(datai[16]), .D1(N309), .S(state), .Y(N7027) );
  mx2a1 U2946 ( .D0(datai[15]), .D1(N308), .S(state), .Y(N7025) );
  mx2a1 U2947 ( .D0(datai[14]), .D1(N307), .S(state), .Y(N7023) );
  mx2a1 U2948 ( .D0(datai[13]), .D1(N306), .S(state), .Y(N7021) );
  mx2a1 U2949 ( .D0(datai[12]), .D1(N305), .S(state), .Y(N7019) );
  mx2a1 U2950 ( .D0(datai[11]), .D1(N304), .S(state), .Y(N7017) );
  mx2a1 U2951 ( .D0(datai[10]), .D1(N303), .S(state), .Y(N7015) );
  mx2a1 U2952 ( .D0(datai[9]), .D1(N302), .S(state), .Y(N7013) );
  mx2a1 U2953 ( .D0(datai[8]), .D1(N301), .S(state), .Y(N7011) );
  mx2a1 U2954 ( .D0(datai[7]), .D1(N300), .S(state), .Y(N7009) );
  mx2a1 U2955 ( .D0(datai[6]), .D1(N299), .S(state), .Y(N7007) );
  mx2a1 U2956 ( .D0(datai[5]), .D1(N298), .S(state), .Y(N7005) );
  mx2a1 U2957 ( .D0(datai[4]), .D1(N297), .S(state), .Y(N7003) );
  mx2a1 U2958 ( .D0(datai[3]), .D1(N296), .S(state), .Y(N7001) );
  mx2a1 U2959 ( .D0(datai[2]), .D1(N295), .S(state), .Y(N6999) );
  mx2a1 U2960 ( .D0(datai[1]), .D1(N294), .S(state), .Y(N6997) );
  mx2a1 U2961 ( .D0(datai[0]), .D1(N293), .S(state), .Y(N6995) );
  ao1f1 U2962 ( .A(n2609), .B(n2462), .C(n2610), .Y(N6993) );
  or4a3 U2963 ( .A(n2611), .B(n2612), .C(n2613), .D(n2614), .Y(N6992) );
  or3a1 U2964 ( .A(n2615), .B(n2616), .C(n2617), .Y(n2614) );
  and2a3 U2965 ( .A(N1354), .B(n2618), .Y(n2617) );
  and2a3 U2966 ( .A(N1334), .B(n2619), .Y(n2616) );
  and2a3 U2967 ( .A(n2620), .B(n201), .Y(n2615) );
  and2a3 U2968 ( .A(reg3[19]), .B(N7058), .Y(n2613) );
  and2a3 U2969 ( .A(n42), .B(n2621), .Y(n2612) );
  and2a3 U2970 ( .A(n2622), .B(N536), .Y(n2611) );
  oa1f1 U2971 ( .A(n2624), .B(n2592), .C(N7058), .Y(n2610) );
  and2a3 U2972 ( .A(n2609), .B(n2625), .Y(n2623) );
  oa1f1 U2973 ( .A(n2626), .B(n2624), .C(n2627), .Y(n2609) );
  or2a1 U2974 ( .A(n2628), .B(n2597), .Y(n2626) );
  or4a3 U2975 ( .A(n2629), .B(n2630), .C(n2631), .D(n2632), .Y(N6990) );
  or3a1 U2976 ( .A(n2633), .B(n2634), .C(n2635), .Y(n2632) );
  and2a3 U2977 ( .A(N1353), .B(n2618), .Y(n2635) );
  and2a3 U2978 ( .A(N1333), .B(n2619), .Y(n2634) );
  and2a3 U2979 ( .A(n2620), .B(n202), .Y(n2633) );
  and2a3 U2980 ( .A(reg3[18]), .B(N7058), .Y(n2631) );
  and2a3 U2981 ( .A(n43), .B(n2621), .Y(n2630) );
  or4a3 U2982 ( .A(n2636), .B(n2637), .C(n2638), .D(n2639), .Y(N6988) );
  or3a1 U2983 ( .A(n2640), .B(n2641), .C(n2642), .Y(n2639) );
  and2a3 U2984 ( .A(N1352), .B(n2618), .Y(n2642) );
  and2a3 U2985 ( .A(N1332), .B(n2619), .Y(n2641) );
  and2a3 U2986 ( .A(n2620), .B(n203), .Y(n2640) );
  and2a3 U2987 ( .A(reg3[17]), .B(N7058), .Y(n2638) );
  and2a3 U2988 ( .A(n44), .B(n2621), .Y(n2637) );
  or4a3 U2989 ( .A(n2643), .B(n2644), .C(n2645), .D(n2646), .Y(N6986) );
  or3a1 U2990 ( .A(n2647), .B(n2648), .C(n2649), .Y(n2646) );
  and2a3 U2991 ( .A(N1351), .B(n2618), .Y(n2649) );
  and2a3 U2992 ( .A(N1331), .B(n2619), .Y(n2648) );
  and2a3 U2993 ( .A(n2620), .B(n204), .Y(n2647) );
  and2a3 U2994 ( .A(reg3[16]), .B(N7058), .Y(n2645) );
  and2a3 U2995 ( .A(n45), .B(n2621), .Y(n2644) );
  or4a3 U2996 ( .A(n2650), .B(n2651), .C(n2652), .D(n2653), .Y(N6984) );
  or3a1 U2997 ( .A(n2654), .B(n2655), .C(n2656), .Y(n2653) );
  and2a3 U2998 ( .A(N1350), .B(n2618), .Y(n2656) );
  and2a3 U2999 ( .A(N1330), .B(n2619), .Y(n2655) );
  and2a3 U3000 ( .A(n2620), .B(n205), .Y(n2654) );
  and2a3 U3001 ( .A(reg3[15]), .B(N7058), .Y(n2652) );
  and2a3 U3002 ( .A(n46), .B(n2621), .Y(n2651) );
  and2a3 U3003 ( .A(n2622), .B(N540), .Y(n2650) );
  or4a3 U3004 ( .A(n2657), .B(n2658), .C(n2659), .D(n2660), .Y(N6982) );
  or3a1 U3005 ( .A(n2661), .B(n2662), .C(n2663), .Y(n2660) );
  and2a3 U3006 ( .A(N1349), .B(n2618), .Y(n2663) );
  and2a3 U3007 ( .A(N1329), .B(n2619), .Y(n2662) );
  and2a3 U3008 ( .A(n2620), .B(n206), .Y(n2661) );
  and2a3 U3009 ( .A(reg3[14]), .B(N7058), .Y(n2659) );
  and2a3 U3010 ( .A(n47), .B(n2621), .Y(n2658) );
  and2a3 U3011 ( .A(n2622), .B(N541), .Y(n2657) );
  or4a3 U3012 ( .A(n2664), .B(n2665), .C(n2666), .D(n2667), .Y(N6980) );
  or3a1 U3013 ( .A(n2668), .B(n2669), .C(n2670), .Y(n2667) );
  and2a3 U3014 ( .A(N1348), .B(n2618), .Y(n2670) );
  and2a3 U3015 ( .A(N1328), .B(n2619), .Y(n2669) );
  and2a3 U3016 ( .A(n2620), .B(n207), .Y(n2668) );
  and2a3 U3017 ( .A(reg3[13]), .B(N7058), .Y(n2666) );
  and2a3 U3018 ( .A(n48), .B(n2621), .Y(n2665) );
  or4a3 U3019 ( .A(n2671), .B(n2672), .C(n2673), .D(n2674), .Y(N6978) );
  or3a1 U3020 ( .A(n2675), .B(n2676), .C(n2677), .Y(n2674) );
  and2a3 U3021 ( .A(N1347), .B(n2618), .Y(n2677) );
  and2a3 U3022 ( .A(N1327), .B(n2619), .Y(n2676) );
  and2a3 U3023 ( .A(n2620), .B(n208), .Y(n2675) );
  and2a3 U3024 ( .A(reg3[12]), .B(N7058), .Y(n2673) );
  and2a3 U3025 ( .A(n49), .B(n2621), .Y(n2672) );
  or4a3 U3026 ( .A(n2678), .B(n2679), .C(n2680), .D(n2681), .Y(N6976) );
  or3a1 U3027 ( .A(n2682), .B(n2683), .C(n2684), .Y(n2681) );
  and2a3 U3028 ( .A(N1346), .B(n2618), .Y(n2684) );
  and2a3 U3029 ( .A(N1326), .B(n2619), .Y(n2683) );
  and2a3 U3030 ( .A(n2620), .B(n209), .Y(n2682) );
  and2a3 U3031 ( .A(reg3[11]), .B(N7058), .Y(n2680) );
  and2a3 U3032 ( .A(n50), .B(n2621), .Y(n2679) );
  and2a3 U3033 ( .A(n2622), .B(N544), .Y(n2678) );
  or4a3 U3034 ( .A(n2685), .B(n2686), .C(n2687), .D(n2688), .Y(N6974) );
  or3a1 U3035 ( .A(n2689), .B(n2690), .C(n2691), .Y(n2688) );
  and2a3 U3036 ( .A(N1345), .B(n2618), .Y(n2691) );
  and2a3 U3037 ( .A(N1325), .B(n2619), .Y(n2690) );
  and2a3 U3038 ( .A(n2620), .B(n210), .Y(n2689) );
  and2a3 U3039 ( .A(reg3[10]), .B(N7058), .Y(n2687) );
  and2a3 U3040 ( .A(n51), .B(n2621), .Y(n2686) );
  and2a3 U3041 ( .A(n2622), .B(N545), .Y(n2685) );
  or4a3 U3042 ( .A(n2692), .B(n2693), .C(n2694), .D(n2695), .Y(N6972) );
  or3a1 U3043 ( .A(n2696), .B(n2697), .C(n2698), .Y(n2695) );
  and2a3 U3044 ( .A(N1344), .B(n2618), .Y(n2698) );
  and2a3 U3045 ( .A(N1324), .B(n2619), .Y(n2697) );
  and2a3 U3046 ( .A(n2620), .B(n211), .Y(n2696) );
  and2a3 U3047 ( .A(reg3[9]), .B(N7058), .Y(n2694) );
  and2a3 U3048 ( .A(n52), .B(n2621), .Y(n2693) );
  or4a3 U3049 ( .A(n2699), .B(n2700), .C(n2701), .D(n2702), .Y(N6970) );
  or3a1 U3050 ( .A(n2703), .B(n2704), .C(n2705), .Y(n2702) );
  and2a3 U3051 ( .A(N1343), .B(n2618), .Y(n2705) );
  and2a3 U3052 ( .A(N1323), .B(n2619), .Y(n2704) );
  and2a3 U3053 ( .A(n2620), .B(n212), .Y(n2703) );
  and2a3 U3054 ( .A(reg3[8]), .B(N7058), .Y(n2701) );
  and2a3 U3055 ( .A(n53), .B(n2621), .Y(n2700) );
  and2a3 U3056 ( .A(n2622), .B(N547), .Y(n2699) );
  or4a3 U3057 ( .A(n2706), .B(n2707), .C(n2708), .D(n2709), .Y(N6968) );
  or3a1 U3058 ( .A(n2710), .B(n2711), .C(n2712), .Y(n2709) );
  and2a3 U3059 ( .A(N1342), .B(n2618), .Y(n2712) );
  and2a3 U3060 ( .A(N1322), .B(n2619), .Y(n2711) );
  and2a3 U3061 ( .A(n2620), .B(n213), .Y(n2710) );
  and2a3 U3062 ( .A(reg3[7]), .B(N7058), .Y(n2708) );
  and2a3 U3063 ( .A(n54), .B(n2621), .Y(n2707) );
  and2a3 U3064 ( .A(n2622), .B(N548), .Y(n2706) );
  or4a3 U3065 ( .A(n2713), .B(n2714), .C(n2715), .D(n2716), .Y(N6966) );
  or3a1 U3066 ( .A(n2717), .B(n2718), .C(n2719), .Y(n2716) );
  and2a3 U3067 ( .A(N1341), .B(n2618), .Y(n2719) );
  and2a3 U3068 ( .A(N1321), .B(n2619), .Y(n2718) );
  and2a3 U3069 ( .A(n2620), .B(n214), .Y(n2717) );
  and2a3 U3070 ( .A(reg3[6]), .B(N7058), .Y(n2715) );
  and2a3 U3071 ( .A(n55), .B(n2621), .Y(n2714) );
  and2a3 U3072 ( .A(n2622), .B(N549), .Y(n2713) );
  or4a3 U3073 ( .A(n2720), .B(n2721), .C(n2722), .D(n2723), .Y(N6964) );
  or3a1 U3074 ( .A(n2724), .B(n2725), .C(n2726), .Y(n2723) );
  and2a3 U3075 ( .A(N1340), .B(n2618), .Y(n2726) );
  and2a3 U3076 ( .A(N1320), .B(n2619), .Y(n2725) );
  and2a3 U3077 ( .A(n2620), .B(n215), .Y(n2724) );
  and2a3 U3078 ( .A(reg3[5]), .B(N7058), .Y(n2722) );
  and2a3 U3079 ( .A(n56), .B(n2621), .Y(n2721) );
  and2a3 U3080 ( .A(n2622), .B(N550), .Y(n2720) );
  or4a3 U3081 ( .A(n2727), .B(n2728), .C(n2729), .D(n2730), .Y(N6962) );
  or4a3 U3082 ( .A(n2731), .B(n2732), .C(n2733), .D(n2734), .Y(n2730) );
  and2a3 U3083 ( .A(N1319), .B(n2619), .Y(n2734) );
  and2a3 U3084 ( .A(n2620), .B(n216), .Y(n2733) );
  and2a3 U3085 ( .A(n2622), .B(N551), .Y(n2732) );
  and2a3 U3086 ( .A(N1339), .B(n2618), .Y(n2731) );
  and2a3 U3087 ( .A(reg3[4]), .B(N7058), .Y(n2729) );
  and2a3 U3088 ( .A(n57), .B(n2621), .Y(n2727) );
  or4a3 U3089 ( .A(n2735), .B(n2736), .C(n2737), .D(n2738), .Y(N6960) );
  or3a1 U3090 ( .A(n2739), .B(n2740), .C(n2741), .Y(n2738) );
  and2a3 U3091 ( .A(N1338), .B(n2618), .Y(n2741) );
  and2a3 U3092 ( .A(N1318), .B(n2619), .Y(n2740) );
  and2a3 U3093 ( .A(n2620), .B(n217), .Y(n2739) );
  and2a3 U3094 ( .A(reg3[3]), .B(N7058), .Y(n2737) );
  and2a3 U3095 ( .A(n58), .B(n2621), .Y(n2736) );
  and2a3 U3096 ( .A(n2622), .B(N552), .Y(n2735) );
  or4a3 U3097 ( .A(n2742), .B(n2728), .C(n2743), .D(n2744), .Y(N6958) );
  or4a3 U3098 ( .A(n2745), .B(n2746), .C(n2747), .D(n2748), .Y(n2744) );
  and2a3 U3099 ( .A(N1317), .B(n2619), .Y(n2748) );
  and2a3 U3100 ( .A(n2620), .B(n218), .Y(n2747) );
  and2a3 U3101 ( .A(N1337), .B(n2618), .Y(n2745) );
  and2a3 U3102 ( .A(reg3[2]), .B(N7058), .Y(n2743) );
  and2a3 U3103 ( .A(N7091), .B(n2749), .Y(n2728) );
  inv1a1 U3104 ( .A(n2750), .Y(n2749) );
  mx2a1 U3105 ( .D0(n2751), .D1(n2752), .S(n2577), .Y(n2750) );
  inv1a1 U3106 ( .A(N555), .Y(n2577) );
  oa1f1 U3107 ( .A(reg2[0]), .B(n2316), .C(n2753), .Y(n2752) );
  and2a3 U3108 ( .A(reg1[0]), .B(n2315), .Y(n2753) );
  and2a3 U3109 ( .A(n2754), .B(n2755), .Y(n2751) );
  mx2a1 U3110 ( .D0(reg2[0]), .D1(reg1[0]), .S(n2756), .Y(n2754) );
  and2a3 U3111 ( .A(n59), .B(n2621), .Y(n2742) );
  or4a3 U3112 ( .A(n2757), .B(n2758), .C(n2759), .D(n2760), .Y(N6956) );
  or3a1 U3113 ( .A(n2761), .B(n2762), .C(n2763), .Y(n2760) );
  and2a3 U3114 ( .A(N1336), .B(n2618), .Y(n2763) );
  and2a3 U3115 ( .A(N1316), .B(n2619), .Y(n2762) );
  and2a3 U3116 ( .A(n2620), .B(n219), .Y(n2761) );
  and2a3 U3117 ( .A(reg3[1]), .B(N7058), .Y(n2759) );
  and2a3 U3118 ( .A(n60), .B(n2621), .Y(n2758) );
  or4a3 U3119 ( .A(n2764), .B(n2765), .C(n2766), .D(n2767), .Y(N6954) );
  or3a1 U3120 ( .A(n2768), .B(n2769), .C(n2770), .Y(n2767) );
  and2a3 U3121 ( .A(N1335), .B(n2618), .Y(n2770) );
  and2a3 U3122 ( .A(N1315), .B(n2619), .Y(n2769) );
  and2a3 U3123 ( .A(n2620), .B(n220), .Y(n2768) );
  and2a3 U3124 ( .A(reg3[0]), .B(N7058), .Y(n2766) );
  and2a3 U3125 ( .A(n61), .B(n2621), .Y(n2765) );
  inv1a1 U3126 ( .A(n2775), .Y(n2774) );
  and3a1 U3127 ( .A(n2589), .B(n2772), .C(n2596), .Y(n2775) );
  and2a3 U3128 ( .A(n2587), .B(n2586), .Y(n2773) );
  or2a1 U3129 ( .A(n2584), .B(n2605), .Y(n2586) );
  inv1a1 U3130 ( .A(n2315), .Y(n2584) );
  or2a1 U3131 ( .A(n2463), .B(n2605), .Y(n2587) );
  inv1a1 U3132 ( .A(n2316), .Y(n2463) );
  inv1a1 U3133 ( .A(n2779), .Y(n2778) );
  or2a1 U3134 ( .A(n2605), .B(N7058), .Y(n2777) );
  ao1f1 U3135 ( .A(n2771), .B(n2628), .C(n2596), .Y(n2776) );
  and2a3 U3136 ( .A(state), .B(n2314), .Y(n2596) );
  or4a3 U3137 ( .A(n2780), .B(n2781), .C(n2782), .D(n2783), .Y(N6920) );
  or3a1 U3138 ( .A(n2784), .B(n2785), .C(n2786), .Y(n2783) );
  and2a3 U3139 ( .A(N584), .B(n2787), .Y(n2786) );
  and2a3 U3140 ( .A(n2788), .B(n192), .Y(n2785) );
  and2a3 U3141 ( .A(n2789), .B(N681), .Y(n2784) );
  and2a3 U3142 ( .A(n33), .B(n2790), .Y(n2782) );
  and2a3 U3143 ( .A(N4683), .B(n2791), .Y(n2781) );
  and2a3 U3144 ( .A(n2792), .B(datai[28]), .Y(n2780) );
  or4a3 U3145 ( .A(n2793), .B(n2794), .C(n2795), .D(n2796), .Y(N6919) );
  or3a1 U3146 ( .A(n2797), .B(n2798), .C(n2799), .Y(n2796) );
  and2a3 U3147 ( .A(N583), .B(n2787), .Y(n2799) );
  and2a3 U3148 ( .A(n2788), .B(n193), .Y(n2798) );
  and2a3 U3149 ( .A(n2789), .B(N680), .Y(n2797) );
  and2a3 U3150 ( .A(n34), .B(n2790), .Y(n2795) );
  and2a3 U3151 ( .A(N4682), .B(n2791), .Y(n2794) );
  and2a3 U3152 ( .A(n2792), .B(datai[27]), .Y(n2793) );
  or4a3 U3153 ( .A(n2800), .B(n2801), .C(n2802), .D(n2803), .Y(N6918) );
  or3a1 U3154 ( .A(n2804), .B(n2805), .C(n2806), .Y(n2803) );
  and2a3 U3155 ( .A(N582), .B(n2787), .Y(n2806) );
  and2a3 U3156 ( .A(n2788), .B(n194), .Y(n2805) );
  and2a3 U3157 ( .A(n2789), .B(N679), .Y(n2804) );
  and2a3 U3158 ( .A(n35), .B(n2790), .Y(n2802) );
  and2a3 U3159 ( .A(N4681), .B(n2791), .Y(n2801) );
  and2a3 U3160 ( .A(n2792), .B(datai[26]), .Y(n2800) );
  or4a3 U3161 ( .A(n2807), .B(n2808), .C(n2809), .D(n2810), .Y(N6917) );
  or3a1 U3162 ( .A(n2811), .B(n2812), .C(n2813), .Y(n2810) );
  and2a3 U3163 ( .A(N581), .B(n2787), .Y(n2813) );
  and2a3 U3164 ( .A(n2788), .B(n195), .Y(n2812) );
  and2a3 U3165 ( .A(n2789), .B(N678), .Y(n2811) );
  and2a3 U3166 ( .A(n36), .B(n2790), .Y(n2809) );
  and2a3 U3167 ( .A(N4680), .B(n2791), .Y(n2808) );
  and2a3 U3168 ( .A(n2792), .B(datai[25]), .Y(n2807) );
  or4a3 U3169 ( .A(n2814), .B(n2815), .C(n2816), .D(n2817), .Y(N6916) );
  or3a1 U3170 ( .A(n2818), .B(n2819), .C(n2820), .Y(n2817) );
  and2a3 U3171 ( .A(N580), .B(n2787), .Y(n2820) );
  and2a3 U3172 ( .A(n2788), .B(n196), .Y(n2819) );
  and2a3 U3173 ( .A(n2789), .B(N677), .Y(n2818) );
  and2a3 U3174 ( .A(n37), .B(n2790), .Y(n2816) );
  and2a3 U3175 ( .A(N4679), .B(n2791), .Y(n2815) );
  and2a3 U3176 ( .A(n2792), .B(datai[24]), .Y(n2814) );
  or4a3 U3177 ( .A(n2821), .B(n2822), .C(n2823), .D(n2824), .Y(N6915) );
  or3a1 U3178 ( .A(n2825), .B(n2826), .C(n2827), .Y(n2824) );
  and2a3 U3179 ( .A(N579), .B(n2787), .Y(n2827) );
  and2a3 U3180 ( .A(n2788), .B(n197), .Y(n2826) );
  and2a3 U3181 ( .A(n2789), .B(N676), .Y(n2825) );
  and2a3 U3182 ( .A(n38), .B(n2790), .Y(n2823) );
  and2a3 U3183 ( .A(N4678), .B(n2791), .Y(n2822) );
  and2a3 U3184 ( .A(n2792), .B(datai[23]), .Y(n2821) );
  or4a3 U3185 ( .A(n2828), .B(n2829), .C(n2830), .D(n2831), .Y(N6914) );
  or3a1 U3186 ( .A(n2832), .B(n2833), .C(n2834), .Y(n2831) );
  and2a3 U3187 ( .A(N578), .B(n2787), .Y(n2834) );
  and2a3 U3188 ( .A(n2788), .B(n198), .Y(n2833) );
  and2a3 U3189 ( .A(n2789), .B(N675), .Y(n2832) );
  and2a3 U3190 ( .A(n39), .B(n2790), .Y(n2830) );
  and2a3 U3191 ( .A(N4677), .B(n2791), .Y(n2829) );
  and2a3 U3192 ( .A(n2792), .B(datai[22]), .Y(n2828) );
  or4a3 U3193 ( .A(n2835), .B(n2836), .C(n2837), .D(n2838), .Y(N6913) );
  or3a1 U3194 ( .A(n2839), .B(n2840), .C(n2841), .Y(n2838) );
  and2a3 U3195 ( .A(N577), .B(n2787), .Y(n2841) );
  and2a3 U3196 ( .A(n2788), .B(n199), .Y(n2840) );
  and2a3 U3197 ( .A(n2789), .B(N674), .Y(n2839) );
  and2a3 U3198 ( .A(n40), .B(n2790), .Y(n2837) );
  and2a3 U3199 ( .A(N4676), .B(n2791), .Y(n2836) );
  and2a3 U3200 ( .A(n2792), .B(datai[21]), .Y(n2835) );
  or4a3 U3201 ( .A(n2842), .B(n2843), .C(n2844), .D(n2845), .Y(N6912) );
  or3a1 U3202 ( .A(n2846), .B(n2847), .C(n2848), .Y(n2845) );
  and2a3 U3203 ( .A(N576), .B(n2787), .Y(n2848) );
  and2a3 U3204 ( .A(n2788), .B(n200), .Y(n2847) );
  and2a3 U3205 ( .A(n2789), .B(N673), .Y(n2846) );
  and2a3 U3206 ( .A(n41), .B(n2790), .Y(n2844) );
  and2a3 U3207 ( .A(N4675), .B(n2791), .Y(n2843) );
  and2a3 U3208 ( .A(n2792), .B(datai[20]), .Y(n2842) );
  ao1f1 U3209 ( .A(n2850), .B(n2851), .C(n2314), .Y(n2849) );
  and2a3 U3210 ( .A(n2597), .B(n2624), .Y(n2851) );
  and2a3 U3211 ( .A(n2627), .B(n2583), .Y(n2850) );
  or4a3 U3212 ( .A(n2852), .B(n2853), .C(n2854), .D(n2855), .Y(N6911) );
  or3a1 U3213 ( .A(n2856), .B(n2857), .C(n2858), .Y(n2855) );
  and2a3 U3214 ( .A(N575), .B(n2787), .Y(n2858) );
  and2a3 U3215 ( .A(n2788), .B(n201), .Y(n2857) );
  and2a3 U3216 ( .A(n2789), .B(N672), .Y(n2856) );
  and2a3 U3217 ( .A(n2790), .B(n42), .Y(n2854) );
  and2a3 U3218 ( .A(N4674), .B(n2791), .Y(n2853) );
  and2a3 U3219 ( .A(n2859), .B(N958), .Y(n2852) );
  or4a3 U3220 ( .A(n2860), .B(n2861), .C(n2862), .D(n2863), .Y(N6910) );
  or3a1 U3221 ( .A(n2864), .B(n2865), .C(n2866), .Y(n2863) );
  and2a3 U3222 ( .A(N574), .B(n2787), .Y(n2866) );
  and2a3 U3223 ( .A(n2788), .B(n202), .Y(n2865) );
  and2a3 U3224 ( .A(n2789), .B(N671), .Y(n2864) );
  and2a3 U3225 ( .A(n2790), .B(n43), .Y(n2862) );
  and2a3 U3226 ( .A(N4673), .B(n2791), .Y(n2861) );
  and2a3 U3227 ( .A(n2859), .B(N957), .Y(n2860) );
  or4a3 U3228 ( .A(n2867), .B(n2868), .C(n2869), .D(n2870), .Y(N6909) );
  or3a1 U3229 ( .A(n2871), .B(n2872), .C(n2873), .Y(n2870) );
  and2a3 U3230 ( .A(N573), .B(n2787), .Y(n2873) );
  and2a3 U3231 ( .A(n2788), .B(n203), .Y(n2872) );
  and2a3 U3232 ( .A(n2789), .B(N670), .Y(n2871) );
  and2a3 U3233 ( .A(n2790), .B(n44), .Y(n2869) );
  and2a3 U3234 ( .A(N4672), .B(n2791), .Y(n2868) );
  and2a3 U3235 ( .A(n2859), .B(N956), .Y(n2867) );
  or4a3 U3236 ( .A(n2874), .B(n2875), .C(n2876), .D(n2877), .Y(N6908) );
  or3a1 U3237 ( .A(n2878), .B(n2879), .C(n2880), .Y(n2877) );
  and2a3 U3238 ( .A(N572), .B(n2787), .Y(n2880) );
  and2a3 U3239 ( .A(n2788), .B(n204), .Y(n2879) );
  and2a3 U3240 ( .A(n2789), .B(N669), .Y(n2878) );
  and2a3 U3241 ( .A(n2790), .B(n45), .Y(n2876) );
  and2a3 U3242 ( .A(N4671), .B(n2791), .Y(n2875) );
  and2a3 U3243 ( .A(n2859), .B(N955), .Y(n2874) );
  or4a3 U3244 ( .A(n2881), .B(n2882), .C(n2883), .D(n2884), .Y(N6907) );
  or3a1 U3245 ( .A(n2885), .B(n2886), .C(n2887), .Y(n2884) );
  and2a3 U3246 ( .A(N571), .B(n2787), .Y(n2887) );
  and2a3 U3247 ( .A(n2788), .B(n205), .Y(n2886) );
  and2a3 U3248 ( .A(n2789), .B(N668), .Y(n2885) );
  and2a3 U3249 ( .A(n2790), .B(n46), .Y(n2883) );
  and2a3 U3250 ( .A(N4670), .B(n2791), .Y(n2882) );
  and2a3 U3251 ( .A(n2859), .B(N954), .Y(n2881) );
  or4a3 U3252 ( .A(n2888), .B(n2889), .C(n2890), .D(n2891), .Y(N6906) );
  or3a1 U3253 ( .A(n2892), .B(n2893), .C(n2894), .Y(n2891) );
  and2a3 U3254 ( .A(N570), .B(n2787), .Y(n2894) );
  and2a3 U3255 ( .A(n2788), .B(n206), .Y(n2893) );
  and2a3 U3256 ( .A(n2789), .B(N667), .Y(n2892) );
  and2a3 U3257 ( .A(n2790), .B(n47), .Y(n2890) );
  and2a3 U3258 ( .A(N4669), .B(n2791), .Y(n2889) );
  and2a3 U3259 ( .A(n2859), .B(N953), .Y(n2888) );
  or4a3 U3260 ( .A(n2895), .B(n2896), .C(n2897), .D(n2898), .Y(N6905) );
  or3a1 U3261 ( .A(n2899), .B(n2900), .C(n2901), .Y(n2898) );
  and2a3 U3262 ( .A(N569), .B(n2787), .Y(n2901) );
  and2a3 U3263 ( .A(n2788), .B(n207), .Y(n2900) );
  and2a3 U3264 ( .A(n2789), .B(N666), .Y(n2899) );
  and2a3 U3265 ( .A(n2790), .B(n48), .Y(n2897) );
  and2a3 U3266 ( .A(N4668), .B(n2791), .Y(n2896) );
  and2a3 U3267 ( .A(n2859), .B(N952), .Y(n2895) );
  or4a3 U3268 ( .A(n2902), .B(n2903), .C(n2904), .D(n2905), .Y(N6904) );
  or3a1 U3269 ( .A(n2906), .B(n2907), .C(n2908), .Y(n2905) );
  and2a3 U3270 ( .A(N568), .B(n2787), .Y(n2908) );
  and2a3 U3271 ( .A(n2788), .B(n208), .Y(n2907) );
  and2a3 U3272 ( .A(n2789), .B(N665), .Y(n2906) );
  and2a3 U3273 ( .A(n2790), .B(n49), .Y(n2904) );
  and2a3 U3274 ( .A(N4667), .B(n2791), .Y(n2903) );
  and2a3 U3275 ( .A(n2859), .B(N951), .Y(n2902) );
  or4a3 U3276 ( .A(n2909), .B(n2910), .C(n2911), .D(n2912), .Y(N6903) );
  or3a1 U3277 ( .A(n2913), .B(n2914), .C(n2915), .Y(n2912) );
  and2a3 U3278 ( .A(N567), .B(n2787), .Y(n2915) );
  and2a3 U3279 ( .A(n2788), .B(n209), .Y(n2914) );
  and2a3 U3280 ( .A(n2789), .B(N664), .Y(n2913) );
  and2a3 U3281 ( .A(n2790), .B(n50), .Y(n2911) );
  and2a3 U3282 ( .A(N4666), .B(n2791), .Y(n2910) );
  and2a3 U3283 ( .A(n2859), .B(N950), .Y(n2909) );
  or4a3 U3284 ( .A(n2916), .B(n2917), .C(n2918), .D(n2919), .Y(N6902) );
  or3a1 U3285 ( .A(n2920), .B(n2921), .C(n2922), .Y(n2919) );
  and2a3 U3286 ( .A(N566), .B(n2787), .Y(n2922) );
  and2a3 U3287 ( .A(n2788), .B(n210), .Y(n2921) );
  and2a3 U3288 ( .A(n2789), .B(N663), .Y(n2920) );
  and2a3 U3289 ( .A(n2790), .B(n51), .Y(n2918) );
  and2a3 U3290 ( .A(N4665), .B(n2791), .Y(n2917) );
  and2a3 U3291 ( .A(n2859), .B(N949), .Y(n2916) );
  or4a3 U3292 ( .A(n2923), .B(n2924), .C(n2925), .D(n2926), .Y(N6901) );
  or3a1 U3293 ( .A(n2927), .B(n2928), .C(n2929), .Y(n2926) );
  and2a3 U3294 ( .A(N565), .B(n2787), .Y(n2929) );
  and2a3 U3295 ( .A(n2788), .B(n211), .Y(n2928) );
  and2a3 U3296 ( .A(n2789), .B(N662), .Y(n2927) );
  and2a3 U3297 ( .A(n2790), .B(n52), .Y(n2925) );
  and2a3 U3298 ( .A(N4664), .B(n2791), .Y(n2924) );
  and2a3 U3299 ( .A(n2859), .B(N948), .Y(n2923) );
  or4a3 U3300 ( .A(n2930), .B(n2931), .C(n2932), .D(n2933), .Y(N6900) );
  or3a1 U3301 ( .A(n2934), .B(n2935), .C(n2936), .Y(n2933) );
  and2a3 U3302 ( .A(N564), .B(n2787), .Y(n2936) );
  and2a3 U3303 ( .A(n2788), .B(n212), .Y(n2935) );
  and2a3 U3304 ( .A(n2789), .B(N661), .Y(n2934) );
  and2a3 U3305 ( .A(n2790), .B(n53), .Y(n2932) );
  and2a3 U3306 ( .A(N4663), .B(n2791), .Y(n2931) );
  and2a3 U3307 ( .A(n2859), .B(N947), .Y(n2930) );
  or4a3 U3308 ( .A(n2937), .B(n2938), .C(n2939), .D(n2940), .Y(N6899) );
  or3a1 U3309 ( .A(n2941), .B(n2942), .C(n2943), .Y(n2940) );
  and2a3 U3310 ( .A(N563), .B(n2787), .Y(n2943) );
  and2a3 U3311 ( .A(n2788), .B(n213), .Y(n2942) );
  and2a3 U3312 ( .A(n2789), .B(N660), .Y(n2941) );
  and2a3 U3313 ( .A(n2790), .B(n54), .Y(n2939) );
  and2a3 U3314 ( .A(N4662), .B(n2791), .Y(n2938) );
  and2a3 U3315 ( .A(n2859), .B(N946), .Y(n2937) );
  or4a3 U3316 ( .A(n2944), .B(n2945), .C(n2946), .D(n2947), .Y(N6898) );
  or3a1 U3317 ( .A(n2948), .B(n2949), .C(n2950), .Y(n2947) );
  and2a3 U3318 ( .A(N562), .B(n2787), .Y(n2950) );
  and2a3 U3319 ( .A(n2788), .B(n214), .Y(n2949) );
  and2a3 U3320 ( .A(n2789), .B(N659), .Y(n2948) );
  and2a3 U3321 ( .A(n2790), .B(n55), .Y(n2946) );
  and2a3 U3322 ( .A(N4661), .B(n2791), .Y(n2945) );
  and2a3 U3323 ( .A(n2859), .B(N945), .Y(n2944) );
  or4a3 U3324 ( .A(n2951), .B(n2952), .C(n2953), .D(n2954), .Y(N6897) );
  or3a1 U3325 ( .A(n2955), .B(n2956), .C(n2957), .Y(n2954) );
  and2a3 U3326 ( .A(N561), .B(n2787), .Y(n2957) );
  and2a3 U3327 ( .A(n2788), .B(n215), .Y(n2956) );
  and2a3 U3328 ( .A(n2789), .B(N658), .Y(n2955) );
  and2a3 U3329 ( .A(n2790), .B(n56), .Y(n2953) );
  and2a3 U3330 ( .A(N4660), .B(n2791), .Y(n2952) );
  and2a3 U3331 ( .A(n2859), .B(N944), .Y(n2951) );
  or4a3 U3332 ( .A(n2958), .B(n2959), .C(n2960), .D(n2961), .Y(N6896) );
  or3a1 U3333 ( .A(n2962), .B(n2963), .C(n2964), .Y(n2961) );
  and2a3 U3334 ( .A(N560), .B(n2787), .Y(n2964) );
  and2a3 U3335 ( .A(n2788), .B(n216), .Y(n2963) );
  and2a3 U3336 ( .A(n2789), .B(N657), .Y(n2962) );
  and2a3 U3337 ( .A(n2790), .B(n57), .Y(n2960) );
  and2a3 U3338 ( .A(N4659), .B(n2791), .Y(n2959) );
  and2a3 U3339 ( .A(n2859), .B(N943), .Y(n2958) );
  or4a3 U3340 ( .A(n2965), .B(n2966), .C(n2967), .D(n2968), .Y(N6895) );
  or3a1 U3341 ( .A(n2969), .B(n2970), .C(n2971), .Y(n2968) );
  and2a3 U3342 ( .A(N559), .B(n2787), .Y(n2971) );
  and2a3 U3343 ( .A(n2788), .B(n217), .Y(n2970) );
  and2a3 U3344 ( .A(n2789), .B(N656), .Y(n2969) );
  and2a3 U3345 ( .A(n2790), .B(n58), .Y(n2967) );
  and2a3 U3346 ( .A(N4658), .B(n2791), .Y(n2966) );
  and2a3 U3347 ( .A(n2859), .B(N942), .Y(n2965) );
  or4a3 U3348 ( .A(n2972), .B(n2973), .C(n2974), .D(n2975), .Y(N6894) );
  or3a1 U3349 ( .A(n2976), .B(n2977), .C(n2978), .Y(n2975) );
  and2a3 U3350 ( .A(N558), .B(n2787), .Y(n2978) );
  and2a3 U3351 ( .A(n2788), .B(n218), .Y(n2977) );
  and2a3 U3352 ( .A(n2789), .B(N655), .Y(n2976) );
  and2a3 U3353 ( .A(n2790), .B(n59), .Y(n2974) );
  and2a3 U3354 ( .A(N4657), .B(n2791), .Y(n2973) );
  and2a3 U3355 ( .A(n2859), .B(N941), .Y(n2972) );
  or4a3 U3356 ( .A(n2979), .B(n2980), .C(n2981), .D(n2982), .Y(N6893) );
  or3a1 U3357 ( .A(n2983), .B(n2984), .C(n2985), .Y(n2982) );
  and2a3 U3358 ( .A(N557), .B(n2787), .Y(n2985) );
  and2a3 U3359 ( .A(n2788), .B(n219), .Y(n2984) );
  and2a3 U3360 ( .A(n2789), .B(N654), .Y(n2983) );
  and2a3 U3361 ( .A(n2790), .B(n60), .Y(n2981) );
  and2a3 U3362 ( .A(N4656), .B(n2791), .Y(n2980) );
  and2a3 U3363 ( .A(n2859), .B(N940), .Y(n2979) );
  or4a3 U3364 ( .A(n2987), .B(n2988), .C(n2989), .D(n2990), .Y(N6892) );
  ao1a1 U3365 ( .A(n220), .B(n2788), .C(n2991), .Y(n2990) );
  and2a3 U3366 ( .A(n2787), .B(N556), .Y(n2991) );
  inv1a1 U3367 ( .A(n2314), .Y(n2462) );
  and2a3 U3368 ( .A(n2604), .B(n2994), .Y(n2993) );
  inv1a1 U3369 ( .A(n2583), .Y(n2994) );
  or3a1 U3370 ( .A(n2995), .B(n2996), .C(n2628), .Y(n2604) );
  or2a1 U3371 ( .A(n2589), .B(n2313), .Y(n2628) );
  or3a1 U3372 ( .A(n2997), .B(n2998), .C(n2999), .Y(n2313) );
  or3a1 U3373 ( .A(n2593), .B(n3000), .C(n3001), .Y(n2589) );
  and3a1 U3374 ( .A(n3002), .B(n3003), .C(n3004), .Y(n2992) );
  and2a3 U3375 ( .A(n2995), .B(n2583), .Y(n2986) );
  and2a3 U3376 ( .A(n2790), .B(n61), .Y(n2989) );
  or4a3 U3377 ( .A(n2581), .B(n2582), .C(n2532), .D(n2580), .Y(n2999) );
  and2a3 U3378 ( .A(N4655), .B(n2791), .Y(n2988) );
  ao1f1 U3379 ( .A(n3000), .B(n2593), .C(n2583), .Y(n3007) );
  or3a1 U3380 ( .A(n2998), .B(n2997), .C(n3001), .Y(n3006) );
  and2a3 U3381 ( .A(n2859), .B(N939), .Y(n2987) );
  and2a3 U3382 ( .A(n2314), .B(n3008), .Y(n2859) );
  inv1a1 U3383 ( .A(n3009), .Y(n3008) );
  ao1f1 U3384 ( .A(n2583), .B(n2597), .C(n2771), .Y(n3009) );
  or2a1 U3385 ( .A(n2597), .B(n2996), .Y(n2771) );
  and2a3 U3386 ( .A(n2602), .B(n2600), .Y(n2583) );
  mx2a1 U3387 ( .D0(d[1]), .D1(N849), .S(n2608), .Y(n2600) );
  xor2a1 U3388 ( .A(n3010), .B(n3011), .Y(N849) );
  mx2a1 U3389 ( .D0(d[0]), .D1(N847), .S(n2608), .Y(n2602) );
  ao1f1 U3390 ( .A(n3010), .B(n3012), .C(n3011), .Y(n2608) );
  xor2a1 U3391 ( .A(n3013), .B(n3014), .Y(n3012) );
  mx2a1 U3392 ( .D0(n3014), .D1(n3015), .S(n3011), .Y(N847) );
  inv1a1 U3393 ( .A(n3010), .Y(n3015) );
  and2a3 U3394 ( .A(n2625), .B(n2605), .Y(n2314) );
  inv1a1 U3395 ( .A(n2607), .Y(n2625) );
  and3a1 U3396 ( .A(n3014), .B(n3010), .C(n3011), .Y(n2607) );
  xor2a1 U3397 ( .A(n3016), .B(n3017), .Y(n3011) );
  and2a3 U3398 ( .A(n3018), .B(n3019), .Y(n3017) );
  xor2a1 U3399 ( .A(n3018), .B(n3019), .Y(n3010) );
  and2a3 U3400 ( .A(n3020), .B(n3021), .Y(n3018) );
  xor2a1 U3401 ( .A(n3021), .B(n3020), .Y(n3014) );
  mx2a1 U3402 ( .D0(N6717), .D1(n3022), .S(n2592), .Y(N6754) );
  inv1a1 U3403 ( .A(n2605), .Y(n2592) );
  oa1f1 U3404 ( .A(n3025), .B(n3026), .C(n3027), .Y(n3024) );
  or4a3 U3405 ( .A(n3028), .B(n3029), .C(n3030), .D(n3031), .Y(n3022) );
  ao1f1 U3406 ( .A(N6305), .B(n3032), .C(n3033), .Y(n3031) );
  ao1f1 U3407 ( .A(n3000), .B(n2590), .C(B), .Y(n3033) );
  or2a1 U3408 ( .A(n3034), .B(n3035), .Y(n2590) );
  inv1a1 U3409 ( .A(n3036), .Y(n3032) );
  oa1f1 U3410 ( .A(n3037), .B(n3038), .C(n3002), .Y(n3030) );
  ao1f1 U3411 ( .A(n3039), .B(n3040), .C(n3041), .Y(n3038) );
  and2a3 U3412 ( .A(n3042), .B(n3043), .Y(n3039) );
  inv1a1 U3413 ( .A(n3044), .Y(n3042) );
  or2a1 U3414 ( .A(n3003), .B(n3045), .Y(n3037) );
  inv1a1 U3415 ( .A(n3046), .Y(n3003) );
  mx2a1 U3416 ( .D0(n3047), .D1(n3048), .S(N6717), .Y(n3029) );
  or2a1 U3417 ( .A(n3034), .B(n2581), .Y(n3048) );
  and3a1 U3418 ( .A(n3004), .B(n3041), .C(n3049), .Y(n3034) );
  or2a1 U3419 ( .A(n3035), .B(n2593), .Y(n3047) );
  and3a1 U3420 ( .A(n3050), .B(n3004), .C(n3049), .Y(n3035) );
  mx2a1 U3421 ( .D0(n3051), .D1(n3052), .S(n3053), .Y(n3028) );
  or3a1 U3422 ( .A(n3054), .B(n3055), .C(n3040), .Y(n3052) );
  and2a3 U3423 ( .A(B), .B(n3004), .Y(n3040) );
  and2a3 U3424 ( .A(n3056), .B(n3045), .Y(n3055) );
  inv1a1 U3425 ( .A(N6175), .Y(n3045) );
  and3a1 U3426 ( .A(n3002), .B(n3050), .C(N6305), .Y(n3054) );
  and2a3 U3427 ( .A(n3056), .B(n3044), .Y(n3051) );
  or4a3 U3428 ( .A(n3057), .B(n3058), .C(n3059), .D(n3060), .Y(n3044) );
  or4a3 U3429 ( .A(n3061), .B(n3062), .C(n3063), .D(n3064), .Y(n3060) );
  or4a3 U3430 ( .A(n3065), .B(n3066), .C(n3067), .D(n3068), .Y(n3064) );
  xor2a1 U3431 ( .A(n2392), .B(n2391), .Y(n3068) );
  xor2a1 U3432 ( .A(n2389), .B(n2388), .Y(n3067) );
  xor2a1 U3433 ( .A(n2323), .B(n2321), .Y(n3066) );
  xor2a1 U3434 ( .A(n2318), .B(n2394), .Y(n3065) );
  or4a3 U3435 ( .A(n3069), .B(n3070), .C(n3071), .D(n3072), .Y(n3063) );
  xor2a1 U3436 ( .A(n2380), .B(n2379), .Y(n3072) );
  xor2a1 U3437 ( .A(n2377), .B(n2376), .Y(n3071) );
  xor2a1 U3438 ( .A(n2386), .B(n2385), .Y(n3070) );
  xor2a1 U3439 ( .A(n2383), .B(n2382), .Y(n3069) );
  or4a3 U3440 ( .A(n3073), .B(n3074), .C(n3075), .D(n3076), .Y(n3062) );
  xor2a1 U3441 ( .A(n2362), .B(n2341), .Y(n3076) );
  xor2a1 U3442 ( .A(n2339), .B(n2337), .Y(n3075) );
  xor2a1 U3443 ( .A(N939), .B(N654), .Y(n3074) );
  xor2a1 U3444 ( .A(n2395), .B(n2364), .Y(n3073) );
  or4a3 U3445 ( .A(n3077), .B(n3078), .C(n3079), .D(n3080), .Y(n3061) );
  xor2a1 U3446 ( .A(n2329), .B(n2328), .Y(n3080) );
  xor2a1 U3447 ( .A(n2326), .B(n2325), .Y(n3079) );
  xor2a1 U3448 ( .A(n2335), .B(n2334), .Y(n3078) );
  xor2a1 U3449 ( .A(n2332), .B(n2331), .Y(n3077) );
  or4a3 U3450 ( .A(n3081), .B(n3082), .C(n3083), .D(n3084), .Y(n3059) );
  or4a3 U3451 ( .A(n3085), .B(n3086), .C(n3087), .D(n3088), .Y(n3084) );
  xor2a1 U3452 ( .A(n2348), .B(n2261), .Y(n3088) );
  inv1a1 U3453 ( .A(N965), .Y(n2348) );
  and2a3 U3454 ( .A(n2624), .B(datai[26]), .Y(N965) );
  xor2a1 U3455 ( .A(n2346), .B(n2259), .Y(n3087) );
  inv1a1 U3456 ( .A(N966), .Y(n2346) );
  and2a3 U3457 ( .A(n2624), .B(datai[27]), .Y(N966) );
  xor2a1 U3458 ( .A(n2352), .B(n2265), .Y(n3086) );
  inv1a1 U3459 ( .A(N963), .Y(n2352) );
  and2a3 U3460 ( .A(n2624), .B(datai[24]), .Y(N963) );
  xor2a1 U3461 ( .A(n2350), .B(n2263), .Y(n3085) );
  inv1a1 U3462 ( .A(N964), .Y(n2350) );
  and2a3 U3463 ( .A(n2624), .B(datai[25]), .Y(N964) );
  or2a1 U3464 ( .A(n3089), .B(n3090), .Y(n3083) );
  xor2a1 U3465 ( .A(n2344), .B(n2257), .Y(n3090) );
  inv1a1 U3466 ( .A(N967), .Y(n2344) );
  and2a3 U3467 ( .A(n2624), .B(datai[28]), .Y(N967) );
  xor2a1 U3468 ( .A(n2342), .B(n2254), .Y(n3089) );
  inv1a1 U3469 ( .A(N683), .Y(n2254) );
  or4a3 U3470 ( .A(n3091), .B(n3092), .C(n3093), .D(n3094), .Y(N683) );
  and2a3 U3471 ( .A(reg1[29]), .B(n3095), .Y(n3094) );
  and2a3 U3472 ( .A(N585), .B(n3096), .Y(n3093) );
  and2a3 U3473 ( .A(reg2[29]), .B(n3097), .Y(n3092) );
  and2a3 U3474 ( .A(reg0[29]), .B(n3098), .Y(n3091) );
  inv1a1 U3475 ( .A(N968), .Y(n2342) );
  and2a3 U3476 ( .A(n2624), .B(datai[29]), .Y(N968) );
  xor2a1 U3477 ( .A(N970), .B(N685), .Y(n3082) );
  and2a3 U3478 ( .A(reg0[31]), .B(n3098), .Y(n3101) );
  and2a3 U3479 ( .A(reg1[31]), .B(n3095), .Y(n3100) );
  and2a3 U3480 ( .A(reg2[31]), .B(n3097), .Y(n3099) );
  and2a3 U3481 ( .A(n2624), .B(datai[31]), .Y(N970) );
  xor2a1 U3482 ( .A(N969), .B(N684), .Y(n3081) );
  and2a3 U3483 ( .A(reg0[30]), .B(n3098), .Y(n3104) );
  and2a3 U3484 ( .A(reg1[30]), .B(n3095), .Y(n3103) );
  and2a3 U3485 ( .A(reg2[30]), .B(n3097), .Y(n3102) );
  and2a3 U3486 ( .A(n2624), .B(datai[30]), .Y(N969) );
  or4a3 U3487 ( .A(n3105), .B(n3106), .C(n3107), .D(n3108), .Y(n3058) );
  xor2a1 U3488 ( .A(n2368), .B(n2367), .Y(n3108) );
  xor2a1 U3489 ( .A(n2365), .B(n2278), .Y(n3107) );
  xor2a1 U3490 ( .A(n2374), .B(n2373), .Y(n3106) );
  xor2a1 U3491 ( .A(n2371), .B(n2370), .Y(n3105) );
  or4a3 U3492 ( .A(n3109), .B(n3110), .C(n3111), .D(n3112), .Y(n3057) );
  xor2a1 U3493 ( .A(n2356), .B(n2269), .Y(n3112) );
  inv1a1 U3494 ( .A(N961), .Y(n2356) );
  and2a3 U3495 ( .A(n2624), .B(datai[22]), .Y(N961) );
  xor2a1 U3496 ( .A(n2354), .B(n2267), .Y(n3111) );
  inv1a1 U3497 ( .A(N962), .Y(n2354) );
  and2a3 U3498 ( .A(n2624), .B(datai[23]), .Y(N962) );
  xor2a1 U3499 ( .A(n2360), .B(n2273), .Y(n3110) );
  inv1a1 U3500 ( .A(N959), .Y(n2360) );
  and2a3 U3501 ( .A(n2624), .B(datai[20]), .Y(N959) );
  xor2a1 U3502 ( .A(n2358), .B(n2271), .Y(n3109) );
  inv1a1 U3503 ( .A(N960), .Y(n2358) );
  and2a3 U3504 ( .A(n2624), .B(datai[21]), .Y(N960) );
  ao1a1 U3505 ( .A(N585), .B(n2597), .C(N5712), .Y(N5776) );
  ao1a1 U3506 ( .A(N584), .B(n2597), .C(N5710), .Y(N5774) );
  ao1a1 U3507 ( .A(N583), .B(n2597), .C(N5708), .Y(N5772) );
  ao1a1 U3508 ( .A(N582), .B(n2597), .C(N5706), .Y(N5770) );
  ao1a1 U3509 ( .A(N581), .B(n2597), .C(N5704), .Y(N5768) );
  ao1a1 U3510 ( .A(N580), .B(n2597), .C(N5702), .Y(N5766) );
  ao1a1 U3511 ( .A(N579), .B(n2597), .C(N5700), .Y(N5764) );
  ao1a1 U3512 ( .A(N578), .B(n2597), .C(N5698), .Y(N5762) );
  ao1a1 U3513 ( .A(N577), .B(n2597), .C(N5696), .Y(N5760) );
  ao1a1 U3514 ( .A(N576), .B(n2597), .C(N5694), .Y(N5758) );
  ao1a1 U3515 ( .A(N575), .B(n2597), .C(N5692), .Y(N5756) );
  ao1a1 U3516 ( .A(N574), .B(n2597), .C(N5690), .Y(N5754) );
  ao1a1 U3517 ( .A(N573), .B(n2597), .C(N5688), .Y(N5752) );
  ao1a1 U3518 ( .A(N572), .B(n2597), .C(N5686), .Y(N5750) );
  ao1a1 U3519 ( .A(N571), .B(n2597), .C(N5684), .Y(N5748) );
  ao1a1 U3520 ( .A(N570), .B(n2597), .C(N5682), .Y(N5746) );
  ao1a1 U3521 ( .A(N569), .B(n2597), .C(N5680), .Y(N5744) );
  ao1a1 U3522 ( .A(N568), .B(n2597), .C(N5678), .Y(N5742) );
  ao1a1 U3523 ( .A(N567), .B(n2597), .C(N5676), .Y(N5740) );
  ao1a1 U3524 ( .A(N566), .B(n2597), .C(N5674), .Y(N5738) );
  ao1a1 U3525 ( .A(N565), .B(n2597), .C(N5672), .Y(N5736) );
  ao1a1 U3526 ( .A(N564), .B(n2597), .C(N5670), .Y(N5734) );
  ao1a1 U3527 ( .A(N563), .B(n2597), .C(N5668), .Y(N5732) );
  ao1a1 U3528 ( .A(N562), .B(n2597), .C(N5666), .Y(N5730) );
  ao1a1 U3529 ( .A(N561), .B(n2597), .C(N5664), .Y(N5728) );
  ao1a1 U3530 ( .A(N560), .B(n2597), .C(N5662), .Y(N5726) );
  ao1a1 U3531 ( .A(N559), .B(n2597), .C(N5660), .Y(N5724) );
  ao1a1 U3532 ( .A(N558), .B(n2597), .C(N5658), .Y(N5722) );
  ao1a1 U3533 ( .A(N557), .B(n2597), .C(N5656), .Y(N5720) );
  ao1a1 U3534 ( .A(N556), .B(n2597), .C(N5654), .Y(N5718) );
  or3a1 U3535 ( .A(n3114), .B(n3115), .C(n3116), .Y(N5780) );
  and2a3 U3536 ( .A(N1059), .B(n2532), .Y(n3116) );
  and2a3 U3537 ( .A(n2627), .B(datai[31]), .Y(n3115) );
  and2a3 U3538 ( .A(n3117), .B(n189), .Y(n3114) );
  or3a1 U3539 ( .A(n3118), .B(n3119), .C(n3120), .Y(N5778) );
  and2a3 U3540 ( .A(N1058), .B(n2532), .Y(n3120) );
  and2a3 U3541 ( .A(n2627), .B(datai[30]), .Y(n3119) );
  and2a3 U3542 ( .A(n3117), .B(n190), .Y(n3118) );
  inv1a1 U3543 ( .A(n3121), .Y(n3117) );
  or4a3 U3544 ( .A(n3122), .B(n3123), .C(n3124), .D(n3125), .Y(N5712) );
  or4a3 U3545 ( .A(n3126), .B(n3127), .C(n3128), .D(n3129), .Y(n3125) );
  or3a1 U3546 ( .A(n3130), .B(n3131), .C(n3132), .Y(n3129) );
  and2a3 U3547 ( .A(N1057), .B(n2532), .Y(n3132) );
  and2a3 U3548 ( .A(N2146), .B(n2998), .Y(n3131) );
  and2a3 U3549 ( .A(N3370), .B(n2593), .Y(n3130) );
  and2a3 U3550 ( .A(N2554), .B(n2580), .Y(n3128) );
  and2a3 U3551 ( .A(N3778), .B(n2997), .Y(n3127) );
  and2a3 U3552 ( .A(N2962), .B(n2581), .Y(n3126) );
  or3a1 U3553 ( .A(n3133), .B(n3134), .C(n3135), .Y(n3124) );
  and2a3 U3554 ( .A(N4186), .B(n2582), .Y(n3135) );
  and2a3 U3555 ( .A(N5002), .B(n3000), .Y(n3134) );
  and2a3 U3556 ( .A(N4594), .B(n3001), .Y(n3133) );
  ao1f1 U3557 ( .A(n2416), .B(n3121), .C(n3136), .Y(n3123) );
  or2a1 U3558 ( .A(n2257), .B(n3137), .Y(n3136) );
  and2a3 U3559 ( .A(reg1[28]), .B(n3095), .Y(n3141) );
  and2a3 U3560 ( .A(N584), .B(n3096), .Y(n3140) );
  and2a3 U3561 ( .A(reg2[28]), .B(n3097), .Y(n3139) );
  and2a3 U3562 ( .A(reg0[28]), .B(n3098), .Y(n3138) );
  ao1f1 U3563 ( .A(n3142), .B(n3143), .C(n2995), .Y(n3121) );
  and2a3 U3564 ( .A(n2779), .B(n3013), .Y(n3142) );
  inv1a1 U3565 ( .A(B), .Y(n3013) );
  inv1a1 U3566 ( .A(n191), .Y(n2416) );
  and2a3 U3567 ( .A(n2627), .B(datai[29]), .Y(n3122) );
  or4a3 U3568 ( .A(n3144), .B(n3145), .C(n3146), .D(n3147), .Y(N5710) );
  or4a3 U3569 ( .A(n3148), .B(n3149), .C(n3150), .D(n3151), .Y(n3147) );
  or3a1 U3570 ( .A(n3152), .B(n3153), .C(n3154), .Y(n3151) );
  and2a3 U3571 ( .A(N1056), .B(n2532), .Y(n3154) );
  and2a3 U3572 ( .A(N2145), .B(n2998), .Y(n3153) );
  and2a3 U3573 ( .A(N3369), .B(n2593), .Y(n3152) );
  and2a3 U3574 ( .A(N2553), .B(n2580), .Y(n3150) );
  and2a3 U3575 ( .A(N3777), .B(n2997), .Y(n3149) );
  and2a3 U3576 ( .A(N2961), .B(n2581), .Y(n3148) );
  or3a1 U3577 ( .A(n3155), .B(n3156), .C(n3157), .Y(n3146) );
  and2a3 U3578 ( .A(N4185), .B(n2582), .Y(n3157) );
  and2a3 U3579 ( .A(N5001), .B(n3000), .Y(n3156) );
  and2a3 U3580 ( .A(N4593), .B(n3001), .Y(n3155) );
  ao1f1 U3581 ( .A(n2259), .B(n3137), .C(n3158), .Y(n3145) );
  or2a1 U3582 ( .A(n3159), .B(n2418), .Y(n3158) );
  inv1a1 U3583 ( .A(n192), .Y(n2418) );
  and2a3 U3584 ( .A(reg1[27]), .B(n3095), .Y(n3163) );
  and2a3 U3585 ( .A(N583), .B(n3096), .Y(n3162) );
  and2a3 U3586 ( .A(reg2[27]), .B(n3097), .Y(n3161) );
  and2a3 U3587 ( .A(reg0[27]), .B(n3098), .Y(n3160) );
  and2a3 U3588 ( .A(n2627), .B(datai[28]), .Y(n3144) );
  or4a3 U3589 ( .A(n3164), .B(n3165), .C(n3166), .D(n3167), .Y(N5708) );
  or4a3 U3590 ( .A(n3168), .B(n3169), .C(n3170), .D(n3171), .Y(n3167) );
  or3a1 U3591 ( .A(n3172), .B(n3173), .C(n3174), .Y(n3171) );
  and2a3 U3592 ( .A(N1055), .B(n2532), .Y(n3174) );
  and2a3 U3593 ( .A(N2144), .B(n2998), .Y(n3173) );
  and2a3 U3594 ( .A(N3368), .B(n2593), .Y(n3172) );
  and2a3 U3595 ( .A(N2552), .B(n2580), .Y(n3170) );
  and2a3 U3596 ( .A(N3776), .B(n2997), .Y(n3169) );
  and2a3 U3597 ( .A(N2960), .B(n2581), .Y(n3168) );
  or3a1 U3598 ( .A(n3175), .B(n3176), .C(n3177), .Y(n3166) );
  and2a3 U3599 ( .A(N4184), .B(n2582), .Y(n3177) );
  and2a3 U3600 ( .A(N5000), .B(n3000), .Y(n3176) );
  and2a3 U3601 ( .A(N4592), .B(n3001), .Y(n3175) );
  ao1f1 U3602 ( .A(n2261), .B(n3137), .C(n3178), .Y(n3165) );
  or2a1 U3603 ( .A(n3159), .B(n2420), .Y(n3178) );
  inv1a1 U3604 ( .A(n193), .Y(n2420) );
  and2a3 U3605 ( .A(reg1[26]), .B(n3095), .Y(n3182) );
  and2a3 U3606 ( .A(N582), .B(n3096), .Y(n3181) );
  and2a3 U3607 ( .A(reg2[26]), .B(n3097), .Y(n3180) );
  and2a3 U3608 ( .A(reg0[26]), .B(n3098), .Y(n3179) );
  and2a3 U3609 ( .A(n2627), .B(datai[27]), .Y(n3164) );
  or4a3 U3610 ( .A(n3183), .B(n3184), .C(n3185), .D(n3186), .Y(N5706) );
  or4a3 U3611 ( .A(n3187), .B(n3188), .C(n3189), .D(n3190), .Y(n3186) );
  or3a1 U3612 ( .A(n3191), .B(n3192), .C(n3193), .Y(n3190) );
  and2a3 U3613 ( .A(N1054), .B(n2532), .Y(n3193) );
  and2a3 U3614 ( .A(N2143), .B(n2998), .Y(n3192) );
  and2a3 U3615 ( .A(N3367), .B(n2593), .Y(n3191) );
  and2a3 U3616 ( .A(N2551), .B(n2580), .Y(n3189) );
  and2a3 U3617 ( .A(N3775), .B(n2997), .Y(n3188) );
  and2a3 U3618 ( .A(N2959), .B(n2581), .Y(n3187) );
  or3a1 U3619 ( .A(n3194), .B(n3195), .C(n3196), .Y(n3185) );
  and2a3 U3620 ( .A(N4183), .B(n2582), .Y(n3196) );
  and2a3 U3621 ( .A(N4999), .B(n3000), .Y(n3195) );
  and2a3 U3622 ( .A(N4591), .B(n3001), .Y(n3194) );
  ao1f1 U3623 ( .A(n2263), .B(n3137), .C(n3197), .Y(n3184) );
  or2a1 U3624 ( .A(n3159), .B(n2422), .Y(n3197) );
  inv1a1 U3625 ( .A(n194), .Y(n2422) );
  and2a3 U3626 ( .A(reg1[25]), .B(n3095), .Y(n3201) );
  and2a3 U3627 ( .A(N581), .B(n3096), .Y(n3200) );
  and2a3 U3628 ( .A(reg2[25]), .B(n3097), .Y(n3199) );
  and2a3 U3629 ( .A(reg0[25]), .B(n3098), .Y(n3198) );
  and2a3 U3630 ( .A(n2627), .B(datai[26]), .Y(n3183) );
  or4a3 U3631 ( .A(n3202), .B(n3203), .C(n3204), .D(n3205), .Y(N5704) );
  or4a3 U3632 ( .A(n3206), .B(n3207), .C(n3208), .D(n3209), .Y(n3205) );
  or3a1 U3633 ( .A(n3210), .B(n3211), .C(n3212), .Y(n3209) );
  and2a3 U3634 ( .A(N1053), .B(n2532), .Y(n3212) );
  and2a3 U3635 ( .A(N2142), .B(n2998), .Y(n3211) );
  and2a3 U3636 ( .A(N3366), .B(n2593), .Y(n3210) );
  and2a3 U3637 ( .A(N2550), .B(n2580), .Y(n3208) );
  and2a3 U3638 ( .A(N3774), .B(n2997), .Y(n3207) );
  and2a3 U3639 ( .A(N2958), .B(n2581), .Y(n3206) );
  or3a1 U3640 ( .A(n3213), .B(n3214), .C(n3215), .Y(n3204) );
  and2a3 U3641 ( .A(N4182), .B(n2582), .Y(n3215) );
  and2a3 U3642 ( .A(N4998), .B(n3000), .Y(n3214) );
  and2a3 U3643 ( .A(N4590), .B(n3001), .Y(n3213) );
  ao1f1 U3644 ( .A(n2265), .B(n3137), .C(n3216), .Y(n3203) );
  or2a1 U3645 ( .A(n3159), .B(n2424), .Y(n3216) );
  inv1a1 U3646 ( .A(n195), .Y(n2424) );
  and2a3 U3647 ( .A(reg1[24]), .B(n3095), .Y(n3220) );
  and2a3 U3648 ( .A(N580), .B(n3096), .Y(n3219) );
  and2a3 U3649 ( .A(reg2[24]), .B(n3097), .Y(n3218) );
  and2a3 U3650 ( .A(reg0[24]), .B(n3098), .Y(n3217) );
  and2a3 U3651 ( .A(n2627), .B(datai[25]), .Y(n3202) );
  or4a3 U3652 ( .A(n3221), .B(n3222), .C(n3223), .D(n3224), .Y(N5702) );
  or4a3 U3653 ( .A(n3225), .B(n3226), .C(n3227), .D(n3228), .Y(n3224) );
  or3a1 U3654 ( .A(n3229), .B(n3230), .C(n3231), .Y(n3228) );
  and2a3 U3655 ( .A(N1052), .B(n2532), .Y(n3231) );
  and2a3 U3656 ( .A(N2141), .B(n2998), .Y(n3230) );
  and2a3 U3657 ( .A(N3365), .B(n2593), .Y(n3229) );
  and2a3 U3658 ( .A(N2549), .B(n2580), .Y(n3227) );
  and2a3 U3659 ( .A(N3773), .B(n2997), .Y(n3226) );
  and2a3 U3660 ( .A(N2957), .B(n2581), .Y(n3225) );
  or3a1 U3661 ( .A(n3232), .B(n3233), .C(n3234), .Y(n3223) );
  and2a3 U3662 ( .A(N4181), .B(n2582), .Y(n3234) );
  and2a3 U3663 ( .A(N4997), .B(n3000), .Y(n3233) );
  and2a3 U3664 ( .A(N4589), .B(n3001), .Y(n3232) );
  ao1f1 U3665 ( .A(n2267), .B(n3137), .C(n3235), .Y(n3222) );
  or2a1 U3666 ( .A(n3159), .B(n2426), .Y(n3235) );
  inv1a1 U3667 ( .A(n196), .Y(n2426) );
  and2a3 U3668 ( .A(reg1[23]), .B(n3095), .Y(n3239) );
  and2a3 U3669 ( .A(N579), .B(n3096), .Y(n3238) );
  and2a3 U3670 ( .A(reg2[23]), .B(n3097), .Y(n3237) );
  and2a3 U3671 ( .A(reg0[23]), .B(n3098), .Y(n3236) );
  and2a3 U3672 ( .A(n2627), .B(datai[24]), .Y(n3221) );
  or4a3 U3673 ( .A(n3240), .B(n3241), .C(n3242), .D(n3243), .Y(N5700) );
  or4a3 U3674 ( .A(n3244), .B(n3245), .C(n3246), .D(n3247), .Y(n3243) );
  or3a1 U3675 ( .A(n3248), .B(n3249), .C(n3250), .Y(n3247) );
  and2a3 U3676 ( .A(N1051), .B(n2532), .Y(n3250) );
  and2a3 U3677 ( .A(N2140), .B(n2998), .Y(n3249) );
  and2a3 U3678 ( .A(N3364), .B(n2593), .Y(n3248) );
  and2a3 U3679 ( .A(N2548), .B(n2580), .Y(n3246) );
  and2a3 U3680 ( .A(N3772), .B(n2997), .Y(n3245) );
  and2a3 U3681 ( .A(N2956), .B(n2581), .Y(n3244) );
  or3a1 U3682 ( .A(n3251), .B(n3252), .C(n3253), .Y(n3242) );
  and2a3 U3683 ( .A(N4180), .B(n2582), .Y(n3253) );
  and2a3 U3684 ( .A(N4996), .B(n3000), .Y(n3252) );
  and2a3 U3685 ( .A(N4588), .B(n3001), .Y(n3251) );
  ao1f1 U3686 ( .A(n2269), .B(n3137), .C(n3254), .Y(n3241) );
  or2a1 U3687 ( .A(n3159), .B(n2428), .Y(n3254) );
  inv1a1 U3688 ( .A(n197), .Y(n2428) );
  and2a3 U3689 ( .A(reg1[22]), .B(n3095), .Y(n3258) );
  and2a3 U3690 ( .A(N578), .B(n3096), .Y(n3257) );
  and2a3 U3691 ( .A(reg2[22]), .B(n3097), .Y(n3256) );
  and2a3 U3692 ( .A(reg0[22]), .B(n3098), .Y(n3255) );
  and2a3 U3693 ( .A(n2627), .B(datai[23]), .Y(n3240) );
  or4a3 U3694 ( .A(n3259), .B(n3260), .C(n3261), .D(n3262), .Y(N5698) );
  or4a3 U3695 ( .A(n3263), .B(n3264), .C(n3265), .D(n3266), .Y(n3262) );
  or3a1 U3696 ( .A(n3267), .B(n3268), .C(n3269), .Y(n3266) );
  and2a3 U3697 ( .A(N1050), .B(n2532), .Y(n3269) );
  and2a3 U3698 ( .A(N2139), .B(n2998), .Y(n3268) );
  and2a3 U3699 ( .A(N3363), .B(n2593), .Y(n3267) );
  and2a3 U3700 ( .A(N2547), .B(n2580), .Y(n3265) );
  and2a3 U3701 ( .A(N3771), .B(n2997), .Y(n3264) );
  and2a3 U3702 ( .A(N2955), .B(n2581), .Y(n3263) );
  or3a1 U3703 ( .A(n3270), .B(n3271), .C(n3272), .Y(n3261) );
  and2a3 U3704 ( .A(N4179), .B(n2582), .Y(n3272) );
  and2a3 U3705 ( .A(N4995), .B(n3000), .Y(n3271) );
  and2a3 U3706 ( .A(N4587), .B(n3001), .Y(n3270) );
  ao1f1 U3707 ( .A(n2271), .B(n3137), .C(n3273), .Y(n3260) );
  or2a1 U3708 ( .A(n3159), .B(n2430), .Y(n3273) );
  inv1a1 U3709 ( .A(n198), .Y(n2430) );
  and2a3 U3710 ( .A(reg1[21]), .B(n3095), .Y(n3277) );
  and2a3 U3711 ( .A(N577), .B(n3096), .Y(n3276) );
  and2a3 U3712 ( .A(reg2[21]), .B(n3097), .Y(n3275) );
  and2a3 U3713 ( .A(reg0[21]), .B(n3098), .Y(n3274) );
  and2a3 U3714 ( .A(n2627), .B(datai[22]), .Y(n3259) );
  or4a3 U3715 ( .A(n3278), .B(n3279), .C(n3280), .D(n3281), .Y(N5696) );
  or4a3 U3716 ( .A(n3282), .B(n3283), .C(n3284), .D(n3285), .Y(n3281) );
  or3a1 U3717 ( .A(n3286), .B(n3287), .C(n3288), .Y(n3285) );
  and2a3 U3718 ( .A(N1049), .B(n2532), .Y(n3288) );
  and2a3 U3719 ( .A(N2138), .B(n2998), .Y(n3287) );
  and2a3 U3720 ( .A(N3362), .B(n2593), .Y(n3286) );
  and2a3 U3721 ( .A(N2546), .B(n2580), .Y(n3284) );
  and2a3 U3722 ( .A(N3770), .B(n2997), .Y(n3283) );
  and2a3 U3723 ( .A(N2954), .B(n2581), .Y(n3282) );
  or3a1 U3724 ( .A(n3289), .B(n3290), .C(n3291), .Y(n3280) );
  and2a3 U3725 ( .A(N4178), .B(n2582), .Y(n3291) );
  and2a3 U3726 ( .A(N4994), .B(n3000), .Y(n3290) );
  and2a3 U3727 ( .A(N4586), .B(n3001), .Y(n3289) );
  ao1f1 U3728 ( .A(n2273), .B(n3137), .C(n3292), .Y(n3279) );
  or2a1 U3729 ( .A(n3159), .B(n2432), .Y(n3292) );
  inv1a1 U3730 ( .A(n199), .Y(n2432) );
  and2a3 U3731 ( .A(reg1[20]), .B(n3095), .Y(n3296) );
  and2a3 U3732 ( .A(N576), .B(n3096), .Y(n3295) );
  and2a3 U3733 ( .A(reg2[20]), .B(n3097), .Y(n3294) );
  and2a3 U3734 ( .A(reg0[20]), .B(n3098), .Y(n3293) );
  and2a3 U3735 ( .A(n2627), .B(datai[21]), .Y(n3278) );
  or4a3 U3736 ( .A(n3297), .B(n3298), .C(n3299), .D(n3300), .Y(N5694) );
  or4a3 U3737 ( .A(n3301), .B(n3302), .C(n3303), .D(n3304), .Y(n3300) );
  or3a1 U3738 ( .A(n3305), .B(n3306), .C(n3307), .Y(n3304) );
  and2a3 U3739 ( .A(N1048), .B(n2532), .Y(n3307) );
  and2a3 U3740 ( .A(N2137), .B(n2998), .Y(n3306) );
  and2a3 U3741 ( .A(N3361), .B(n2593), .Y(n3305) );
  and2a3 U3742 ( .A(N2545), .B(n2580), .Y(n3303) );
  and2a3 U3743 ( .A(N3769), .B(n2997), .Y(n3302) );
  and2a3 U3744 ( .A(N2953), .B(n2581), .Y(n3301) );
  or3a1 U3745 ( .A(n3308), .B(n3309), .C(n3310), .Y(n3299) );
  and2a3 U3746 ( .A(N4177), .B(n2582), .Y(n3310) );
  and2a3 U3747 ( .A(N4993), .B(n3000), .Y(n3309) );
  and2a3 U3748 ( .A(N4585), .B(n3001), .Y(n3308) );
  ao1f1 U3749 ( .A(n3159), .B(n2434), .C(n3311), .Y(n3298) );
  or2a1 U3750 ( .A(n2278), .B(n3137), .Y(n3311) );
  and2a3 U3751 ( .A(N575), .B(n3096), .Y(n3315) );
  and2a3 U3752 ( .A(n3097), .B(reg2[19]), .Y(n3314) );
  and2a3 U3753 ( .A(n3095), .B(reg1[19]), .Y(n3313) );
  and2a3 U3754 ( .A(reg0[19]), .B(n3098), .Y(n3312) );
  inv1a1 U3755 ( .A(n200), .Y(n2434) );
  and2a3 U3756 ( .A(n2627), .B(datai[20]), .Y(n3297) );
  and2a3 U3757 ( .A(n2624), .B(n2996), .Y(n2627) );
  or4a3 U3758 ( .A(n3316), .B(n3317), .C(n3318), .D(n3319), .Y(N5692) );
  or4a3 U3759 ( .A(n3320), .B(n3321), .C(n3322), .D(n3323), .Y(n3319) );
  or3a1 U3760 ( .A(n3324), .B(n3325), .C(n3326), .Y(n3323) );
  and2a3 U3761 ( .A(N1047), .B(n2532), .Y(n3326) );
  and2a3 U3762 ( .A(N2136), .B(n2998), .Y(n3325) );
  and2a3 U3763 ( .A(N3360), .B(n2593), .Y(n3324) );
  and2a3 U3764 ( .A(N2544), .B(n2580), .Y(n3322) );
  and2a3 U3765 ( .A(N3768), .B(n2997), .Y(n3321) );
  and2a3 U3766 ( .A(N2952), .B(n2581), .Y(n3320) );
  or3a1 U3767 ( .A(n3327), .B(n3328), .C(n3329), .Y(n3318) );
  and2a3 U3768 ( .A(N4176), .B(n2582), .Y(n3329) );
  and2a3 U3769 ( .A(N4992), .B(n3000), .Y(n3328) );
  and2a3 U3770 ( .A(N4584), .B(n3001), .Y(n3327) );
  ao1f1 U3771 ( .A(n3159), .B(n2438), .C(n3330), .Y(n3317) );
  or2a1 U3772 ( .A(n2367), .B(n3137), .Y(n3330) );
  inv1a1 U3773 ( .A(N672), .Y(n2367) );
  and2a3 U3774 ( .A(N574), .B(n3096), .Y(n3334) );
  and2a3 U3775 ( .A(reg2[18]), .B(n3097), .Y(n3333) );
  and2a3 U3776 ( .A(reg1[18]), .B(n3095), .Y(n3332) );
  and2a3 U3777 ( .A(reg0[18]), .B(n3098), .Y(n3331) );
  inv1a1 U3778 ( .A(n201), .Y(n2438) );
  and2a3 U3779 ( .A(n2996), .B(N958), .Y(n3316) );
  oa1f1 U3780 ( .A(N536), .B(n3143), .C(n3335), .Y(n2365) );
  and2a3 U3781 ( .A(n2624), .B(datai[19]), .Y(n3335) );
  or4a3 U3782 ( .A(n3336), .B(n3337), .C(n3338), .D(n3339), .Y(N5690) );
  or4a3 U3783 ( .A(n3340), .B(n3341), .C(n3342), .D(n3343), .Y(n3339) );
  or3a1 U3784 ( .A(n3344), .B(n3345), .C(n3346), .Y(n3343) );
  and2a3 U3785 ( .A(N1046), .B(n2532), .Y(n3346) );
  and2a3 U3786 ( .A(N2135), .B(n2998), .Y(n3345) );
  and2a3 U3787 ( .A(N3359), .B(n2593), .Y(n3344) );
  and2a3 U3788 ( .A(N2543), .B(n2580), .Y(n3342) );
  and2a3 U3789 ( .A(N3767), .B(n2997), .Y(n3341) );
  and2a3 U3790 ( .A(N2951), .B(n2581), .Y(n3340) );
  or3a1 U3791 ( .A(n3347), .B(n3348), .C(n3349), .Y(n3338) );
  and2a3 U3792 ( .A(N4175), .B(n2582), .Y(n3349) );
  and2a3 U3793 ( .A(N4991), .B(n3000), .Y(n3348) );
  and2a3 U3794 ( .A(N4583), .B(n3001), .Y(n3347) );
  ao1f1 U3795 ( .A(n3159), .B(n2440), .C(n3350), .Y(n3337) );
  or2a1 U3796 ( .A(n2370), .B(n3137), .Y(n3350) );
  inv1a1 U3797 ( .A(N671), .Y(n2370) );
  and2a3 U3798 ( .A(N573), .B(n3096), .Y(n3354) );
  and2a3 U3799 ( .A(reg2[17]), .B(n3097), .Y(n3353) );
  and2a3 U3800 ( .A(reg1[17]), .B(n3095), .Y(n3352) );
  and2a3 U3801 ( .A(reg0[17]), .B(n3098), .Y(n3351) );
  inv1a1 U3802 ( .A(n202), .Y(n2440) );
  and2a3 U3803 ( .A(n2996), .B(N957), .Y(n3336) );
  oa1f1 U3804 ( .A(N537), .B(n3143), .C(n3355), .Y(n2368) );
  and2a3 U3805 ( .A(n2624), .B(datai[18]), .Y(n3355) );
  or4a3 U3806 ( .A(n3356), .B(n3357), .C(n3358), .D(n3359), .Y(N5688) );
  or4a3 U3807 ( .A(n3360), .B(n3361), .C(n3362), .D(n3363), .Y(n3359) );
  or3a1 U3808 ( .A(n3364), .B(n3365), .C(n3366), .Y(n3363) );
  and2a3 U3809 ( .A(N1045), .B(n2532), .Y(n3366) );
  and2a3 U3810 ( .A(N2134), .B(n2998), .Y(n3365) );
  and2a3 U3811 ( .A(N3358), .B(n2593), .Y(n3364) );
  and2a3 U3812 ( .A(N2542), .B(n2580), .Y(n3362) );
  and2a3 U3813 ( .A(N3766), .B(n2997), .Y(n3361) );
  and2a3 U3814 ( .A(N2950), .B(n2581), .Y(n3360) );
  or3a1 U3815 ( .A(n3367), .B(n3368), .C(n3369), .Y(n3358) );
  and2a3 U3816 ( .A(N4174), .B(n2582), .Y(n3369) );
  and2a3 U3817 ( .A(N4990), .B(n3000), .Y(n3368) );
  and2a3 U3818 ( .A(N4582), .B(n3001), .Y(n3367) );
  ao1f1 U3819 ( .A(n3159), .B(n2442), .C(n3370), .Y(n3357) );
  or2a1 U3820 ( .A(n2373), .B(n3137), .Y(n3370) );
  inv1a1 U3821 ( .A(N670), .Y(n2373) );
  and2a3 U3822 ( .A(N572), .B(n3096), .Y(n3374) );
  and2a3 U3823 ( .A(reg2[16]), .B(n3097), .Y(n3373) );
  and2a3 U3824 ( .A(reg1[16]), .B(n3095), .Y(n3372) );
  and2a3 U3825 ( .A(reg0[16]), .B(n3098), .Y(n3371) );
  inv1a1 U3826 ( .A(n203), .Y(n2442) );
  and2a3 U3827 ( .A(n2996), .B(N956), .Y(n3356) );
  oa1f1 U3828 ( .A(N538), .B(n3143), .C(n3375), .Y(n2371) );
  and2a3 U3829 ( .A(n2624), .B(datai[17]), .Y(n3375) );
  or4a3 U3830 ( .A(n3376), .B(n3377), .C(n3378), .D(n3379), .Y(N5686) );
  or4a3 U3831 ( .A(n3380), .B(n3381), .C(n3382), .D(n3383), .Y(n3379) );
  or3a1 U3832 ( .A(n3384), .B(n3385), .C(n3386), .Y(n3383) );
  and2a3 U3833 ( .A(N1044), .B(n2532), .Y(n3386) );
  and2a3 U3834 ( .A(N2133), .B(n2998), .Y(n3385) );
  and2a3 U3835 ( .A(N3357), .B(n2593), .Y(n3384) );
  and2a3 U3836 ( .A(N2541), .B(n2580), .Y(n3382) );
  and2a3 U3837 ( .A(N3765), .B(n2997), .Y(n3381) );
  and2a3 U3838 ( .A(N2949), .B(n2581), .Y(n3380) );
  or3a1 U3839 ( .A(n3387), .B(n3388), .C(n3389), .Y(n3378) );
  and2a3 U3840 ( .A(N4173), .B(n2582), .Y(n3389) );
  and2a3 U3841 ( .A(N4989), .B(n3000), .Y(n3388) );
  and2a3 U3842 ( .A(N4581), .B(n3001), .Y(n3387) );
  ao1f1 U3843 ( .A(n3159), .B(n2444), .C(n3390), .Y(n3377) );
  or2a1 U3844 ( .A(n2376), .B(n3137), .Y(n3390) );
  inv1a1 U3845 ( .A(N669), .Y(n2376) );
  and2a3 U3846 ( .A(N571), .B(n3096), .Y(n3394) );
  and2a3 U3847 ( .A(reg2[15]), .B(n3097), .Y(n3393) );
  and2a3 U3848 ( .A(reg1[15]), .B(n3095), .Y(n3392) );
  and2a3 U3849 ( .A(reg0[15]), .B(n3098), .Y(n3391) );
  inv1a1 U3850 ( .A(n204), .Y(n2444) );
  and2a3 U3851 ( .A(n2996), .B(N955), .Y(n3376) );
  oa1f1 U3852 ( .A(N539), .B(n3143), .C(n3395), .Y(n2374) );
  and2a3 U3853 ( .A(n2624), .B(datai[16]), .Y(n3395) );
  or4a3 U3854 ( .A(n3396), .B(n3397), .C(n3398), .D(n3399), .Y(N5684) );
  or4a3 U3855 ( .A(n3400), .B(n3401), .C(n3402), .D(n3403), .Y(n3399) );
  or3a1 U3856 ( .A(n3404), .B(n3405), .C(n3406), .Y(n3403) );
  and2a3 U3857 ( .A(N1043), .B(n2532), .Y(n3406) );
  and2a3 U3858 ( .A(N2132), .B(n2998), .Y(n3405) );
  and2a3 U3859 ( .A(N3356), .B(n2593), .Y(n3404) );
  and2a3 U3860 ( .A(N2540), .B(n2580), .Y(n3402) );
  and2a3 U3861 ( .A(N3764), .B(n2997), .Y(n3401) );
  and2a3 U3862 ( .A(N2948), .B(n2581), .Y(n3400) );
  or3a1 U3863 ( .A(n3407), .B(n3408), .C(n3409), .Y(n3398) );
  and2a3 U3864 ( .A(N4172), .B(n2582), .Y(n3409) );
  and2a3 U3865 ( .A(N4988), .B(n3000), .Y(n3408) );
  and2a3 U3866 ( .A(N4580), .B(n3001), .Y(n3407) );
  ao1f1 U3867 ( .A(n3159), .B(n2446), .C(n3410), .Y(n3397) );
  or2a1 U3868 ( .A(n2379), .B(n3137), .Y(n3410) );
  inv1a1 U3869 ( .A(N668), .Y(n2379) );
  and2a3 U3870 ( .A(N570), .B(n3096), .Y(n3414) );
  and2a3 U3871 ( .A(reg2[14]), .B(n3097), .Y(n3413) );
  and2a3 U3872 ( .A(reg1[14]), .B(n3095), .Y(n3412) );
  and2a3 U3873 ( .A(reg0[14]), .B(n3098), .Y(n3411) );
  inv1a1 U3874 ( .A(n205), .Y(n2446) );
  and2a3 U3875 ( .A(n2996), .B(N954), .Y(n3396) );
  oa1f1 U3876 ( .A(N540), .B(n3143), .C(n3415), .Y(n2377) );
  and2a3 U3877 ( .A(n2624), .B(datai[15]), .Y(n3415) );
  or4a3 U3878 ( .A(n3416), .B(n3417), .C(n3418), .D(n3419), .Y(N5682) );
  or4a3 U3879 ( .A(n3420), .B(n3421), .C(n3422), .D(n3423), .Y(n3419) );
  or3a1 U3880 ( .A(n3424), .B(n3425), .C(n3426), .Y(n3423) );
  and2a3 U3881 ( .A(N1042), .B(n2532), .Y(n3426) );
  and2a3 U3882 ( .A(N2131), .B(n2998), .Y(n3425) );
  and2a3 U3883 ( .A(N3355), .B(n2593), .Y(n3424) );
  and2a3 U3884 ( .A(N2539), .B(n2580), .Y(n3422) );
  and2a3 U3885 ( .A(N3763), .B(n2997), .Y(n3421) );
  and2a3 U3886 ( .A(N2947), .B(n2581), .Y(n3420) );
  or3a1 U3887 ( .A(n3427), .B(n3428), .C(n3429), .Y(n3418) );
  and2a3 U3888 ( .A(N4171), .B(n2582), .Y(n3429) );
  and2a3 U3889 ( .A(N4987), .B(n3000), .Y(n3428) );
  and2a3 U3890 ( .A(N4579), .B(n3001), .Y(n3427) );
  ao1f1 U3891 ( .A(n3159), .B(n2448), .C(n3430), .Y(n3417) );
  or2a1 U3892 ( .A(n2382), .B(n3137), .Y(n3430) );
  inv1a1 U3893 ( .A(N667), .Y(n2382) );
  and2a3 U3894 ( .A(N569), .B(n3096), .Y(n3434) );
  and2a3 U3895 ( .A(reg2[13]), .B(n3097), .Y(n3433) );
  and2a3 U3896 ( .A(reg1[13]), .B(n3095), .Y(n3432) );
  and2a3 U3897 ( .A(reg0[13]), .B(n3098), .Y(n3431) );
  inv1a1 U3898 ( .A(n206), .Y(n2448) );
  and2a3 U3899 ( .A(n2996), .B(N953), .Y(n3416) );
  oa1f1 U3900 ( .A(N541), .B(n3143), .C(n3435), .Y(n2380) );
  and2a3 U3901 ( .A(n2624), .B(datai[14]), .Y(n3435) );
  or4a3 U3902 ( .A(n3436), .B(n3437), .C(n3438), .D(n3439), .Y(N5680) );
  or4a3 U3903 ( .A(n3440), .B(n3441), .C(n3442), .D(n3443), .Y(n3439) );
  or3a1 U3904 ( .A(n3444), .B(n3445), .C(n3446), .Y(n3443) );
  and2a3 U3905 ( .A(N1041), .B(n2532), .Y(n3446) );
  and2a3 U3906 ( .A(N2130), .B(n2998), .Y(n3445) );
  and2a3 U3907 ( .A(N3354), .B(n2593), .Y(n3444) );
  and2a3 U3908 ( .A(N2538), .B(n2580), .Y(n3442) );
  and2a3 U3909 ( .A(N3762), .B(n2997), .Y(n3441) );
  and2a3 U3910 ( .A(N2946), .B(n2581), .Y(n3440) );
  or3a1 U3911 ( .A(n3447), .B(n3448), .C(n3449), .Y(n3438) );
  and2a3 U3912 ( .A(N4170), .B(n2582), .Y(n3449) );
  and2a3 U3913 ( .A(N4986), .B(n3000), .Y(n3448) );
  and2a3 U3914 ( .A(N4578), .B(n3001), .Y(n3447) );
  ao1f1 U3915 ( .A(n3159), .B(n2450), .C(n3450), .Y(n3437) );
  or2a1 U3916 ( .A(n2385), .B(n3137), .Y(n3450) );
  inv1a1 U3917 ( .A(N666), .Y(n2385) );
  and2a3 U3918 ( .A(N568), .B(n3096), .Y(n3454) );
  and2a3 U3919 ( .A(reg2[12]), .B(n3097), .Y(n3453) );
  and2a3 U3920 ( .A(reg1[12]), .B(n3095), .Y(n3452) );
  and2a3 U3921 ( .A(reg0[12]), .B(n3098), .Y(n3451) );
  inv1a1 U3922 ( .A(n207), .Y(n2450) );
  and2a3 U3923 ( .A(n2996), .B(N952), .Y(n3436) );
  oa1f1 U3924 ( .A(N542), .B(n3143), .C(n3455), .Y(n2383) );
  and2a3 U3925 ( .A(n2624), .B(datai[13]), .Y(n3455) );
  or4a3 U3926 ( .A(n3456), .B(n3457), .C(n3458), .D(n3459), .Y(N5678) );
  or4a3 U3927 ( .A(n3460), .B(n3461), .C(n3462), .D(n3463), .Y(n3459) );
  or3a1 U3928 ( .A(n3464), .B(n3465), .C(n3466), .Y(n3463) );
  and2a3 U3929 ( .A(N1040), .B(n2532), .Y(n3466) );
  and2a3 U3930 ( .A(N2129), .B(n2998), .Y(n3465) );
  and2a3 U3931 ( .A(N3353), .B(n2593), .Y(n3464) );
  and2a3 U3932 ( .A(N2537), .B(n2580), .Y(n3462) );
  and2a3 U3933 ( .A(N3761), .B(n2997), .Y(n3461) );
  and2a3 U3934 ( .A(N2945), .B(n2581), .Y(n3460) );
  or3a1 U3935 ( .A(n3467), .B(n3468), .C(n3469), .Y(n3458) );
  and2a3 U3936 ( .A(N4169), .B(n2582), .Y(n3469) );
  and2a3 U3937 ( .A(N4985), .B(n3000), .Y(n3468) );
  and2a3 U3938 ( .A(N4577), .B(n3001), .Y(n3467) );
  ao1f1 U3939 ( .A(n3159), .B(n2452), .C(n3470), .Y(n3457) );
  or2a1 U3940 ( .A(n2388), .B(n3137), .Y(n3470) );
  inv1a1 U3941 ( .A(N665), .Y(n2388) );
  and2a3 U3942 ( .A(N567), .B(n3096), .Y(n3474) );
  and2a3 U3943 ( .A(reg2[11]), .B(n3097), .Y(n3473) );
  and2a3 U3944 ( .A(reg1[11]), .B(n3095), .Y(n3472) );
  and2a3 U3945 ( .A(reg0[11]), .B(n3098), .Y(n3471) );
  inv1a1 U3946 ( .A(n208), .Y(n2452) );
  and2a3 U3947 ( .A(n2996), .B(N951), .Y(n3456) );
  oa1f1 U3948 ( .A(N543), .B(n3143), .C(n3475), .Y(n2386) );
  and2a3 U3949 ( .A(n2624), .B(datai[12]), .Y(n3475) );
  or4a3 U3950 ( .A(n3476), .B(n3477), .C(n3478), .D(n3479), .Y(N5676) );
  or4a3 U3951 ( .A(n3480), .B(n3481), .C(n3482), .D(n3483), .Y(n3479) );
  or3a1 U3952 ( .A(n3484), .B(n3485), .C(n3486), .Y(n3483) );
  and2a3 U3953 ( .A(N1039), .B(n2532), .Y(n3486) );
  and2a3 U3954 ( .A(N2128), .B(n2998), .Y(n3485) );
  and2a3 U3955 ( .A(N3352), .B(n2593), .Y(n3484) );
  and2a3 U3956 ( .A(N2536), .B(n2580), .Y(n3482) );
  and2a3 U3957 ( .A(N3760), .B(n2997), .Y(n3481) );
  and2a3 U3958 ( .A(N2944), .B(n2581), .Y(n3480) );
  or3a1 U3959 ( .A(n3487), .B(n3488), .C(n3489), .Y(n3478) );
  and2a3 U3960 ( .A(N4168), .B(n2582), .Y(n3489) );
  and2a3 U3961 ( .A(N4984), .B(n3000), .Y(n3488) );
  and2a3 U3962 ( .A(N4576), .B(n3001), .Y(n3487) );
  ao1f1 U3963 ( .A(n3159), .B(n2454), .C(n3490), .Y(n3477) );
  or2a1 U3964 ( .A(n2391), .B(n3137), .Y(n3490) );
  inv1a1 U3965 ( .A(N664), .Y(n2391) );
  and2a3 U3966 ( .A(N566), .B(n3096), .Y(n3494) );
  and2a3 U3967 ( .A(reg2[10]), .B(n3097), .Y(n3493) );
  and2a3 U3968 ( .A(reg1[10]), .B(n3095), .Y(n3492) );
  and2a3 U3969 ( .A(reg0[10]), .B(n3098), .Y(n3491) );
  inv1a1 U3970 ( .A(n209), .Y(n2454) );
  and2a3 U3971 ( .A(n2996), .B(N950), .Y(n3476) );
  oa1f1 U3972 ( .A(N544), .B(n3143), .C(n3495), .Y(n2389) );
  and2a3 U3973 ( .A(n2624), .B(datai[11]), .Y(n3495) );
  or4a3 U3974 ( .A(n3496), .B(n3497), .C(n3498), .D(n3499), .Y(N5674) );
  or4a3 U3975 ( .A(n3500), .B(n3501), .C(n3502), .D(n3503), .Y(n3499) );
  or3a1 U3976 ( .A(n3504), .B(n3505), .C(n3506), .Y(n3503) );
  and2a3 U3977 ( .A(N1038), .B(n2532), .Y(n3506) );
  and2a3 U3978 ( .A(N2127), .B(n2998), .Y(n3505) );
  and2a3 U3979 ( .A(N3351), .B(n2593), .Y(n3504) );
  and2a3 U3980 ( .A(N2535), .B(n2580), .Y(n3502) );
  and2a3 U3981 ( .A(N3759), .B(n2997), .Y(n3501) );
  and2a3 U3982 ( .A(N2943), .B(n2581), .Y(n3500) );
  or3a1 U3983 ( .A(n3507), .B(n3508), .C(n3509), .Y(n3498) );
  and2a3 U3984 ( .A(N4167), .B(n2582), .Y(n3509) );
  and2a3 U3985 ( .A(N4983), .B(n3000), .Y(n3508) );
  and2a3 U3986 ( .A(N4575), .B(n3001), .Y(n3507) );
  ao1f1 U3987 ( .A(n3159), .B(n2456), .C(n3510), .Y(n3497) );
  or2a1 U3988 ( .A(n2394), .B(n3137), .Y(n3510) );
  inv1a1 U3989 ( .A(N663), .Y(n2394) );
  and2a3 U3990 ( .A(N565), .B(n3096), .Y(n3514) );
  and2a3 U3991 ( .A(n3097), .B(reg2[9]), .Y(n3513) );
  and2a3 U3992 ( .A(n3095), .B(reg1[9]), .Y(n3512) );
  and2a3 U3993 ( .A(reg0[9]), .B(n3098), .Y(n3511) );
  inv1a1 U3994 ( .A(n210), .Y(n2456) );
  and2a3 U3995 ( .A(n2996), .B(N949), .Y(n3496) );
  oa1f1 U3996 ( .A(N545), .B(n3143), .C(n3515), .Y(n2392) );
  and2a3 U3997 ( .A(n2624), .B(datai[10]), .Y(n3515) );
  or4a3 U3998 ( .A(n3516), .B(n3517), .C(n3518), .D(n3519), .Y(N5672) );
  or4a3 U3999 ( .A(n3520), .B(n3521), .C(n3522), .D(n3523), .Y(n3519) );
  or3a1 U4000 ( .A(n3524), .B(n3525), .C(n3526), .Y(n3523) );
  and2a3 U4001 ( .A(N1037), .B(n2532), .Y(n3526) );
  and2a3 U4002 ( .A(N2126), .B(n2998), .Y(n3525) );
  and2a3 U4003 ( .A(N3350), .B(n2593), .Y(n3524) );
  and2a3 U4004 ( .A(N2534), .B(n2580), .Y(n3522) );
  and2a3 U4005 ( .A(N3758), .B(n2997), .Y(n3521) );
  and2a3 U4006 ( .A(N2942), .B(n2581), .Y(n3520) );
  or3a1 U4007 ( .A(n3527), .B(n3528), .C(n3529), .Y(n3518) );
  and2a3 U4008 ( .A(N4166), .B(n2582), .Y(n3529) );
  and2a3 U4009 ( .A(N4982), .B(n3000), .Y(n3528) );
  and2a3 U4010 ( .A(N4574), .B(n3001), .Y(n3527) );
  ao1f1 U4011 ( .A(n3159), .B(n2398), .C(n3530), .Y(n3517) );
  or2a1 U4012 ( .A(n2321), .B(n3137), .Y(n3530) );
  inv1a1 U4013 ( .A(N662), .Y(n2321) );
  and2a3 U4014 ( .A(N564), .B(n3096), .Y(n3534) );
  and2a3 U4015 ( .A(n3097), .B(reg2[8]), .Y(n3533) );
  and2a3 U4016 ( .A(n3095), .B(reg1[8]), .Y(n3532) );
  and2a3 U4017 ( .A(reg0[8]), .B(n3098), .Y(n3531) );
  inv1a1 U4018 ( .A(n211), .Y(n2398) );
  and2a3 U4019 ( .A(n2996), .B(N948), .Y(n3516) );
  oa1f1 U4020 ( .A(N546), .B(n3143), .C(n3535), .Y(n2318) );
  and2a3 U4021 ( .A(n2624), .B(datai[9]), .Y(n3535) );
  or4a3 U4022 ( .A(n3536), .B(n3537), .C(n3538), .D(n3539), .Y(N5670) );
  or4a3 U4023 ( .A(n3540), .B(n3541), .C(n3542), .D(n3543), .Y(n3539) );
  or3a1 U4024 ( .A(n3544), .B(n3545), .C(n3546), .Y(n3543) );
  and2a3 U4025 ( .A(N1036), .B(n2532), .Y(n3546) );
  and2a3 U4026 ( .A(N2125), .B(n2998), .Y(n3545) );
  and2a3 U4027 ( .A(N3349), .B(n2593), .Y(n3544) );
  and2a3 U4028 ( .A(N2533), .B(n2580), .Y(n3542) );
  and2a3 U4029 ( .A(N3757), .B(n2997), .Y(n3541) );
  and2a3 U4030 ( .A(N2941), .B(n2581), .Y(n3540) );
  or3a1 U4031 ( .A(n3547), .B(n3548), .C(n3549), .Y(n3538) );
  and2a3 U4032 ( .A(N4165), .B(n2582), .Y(n3549) );
  and2a3 U4033 ( .A(N4981), .B(n3000), .Y(n3548) );
  and2a3 U4034 ( .A(N4573), .B(n3001), .Y(n3547) );
  ao1f1 U4035 ( .A(n3159), .B(n2402), .C(n3550), .Y(n3537) );
  or2a1 U4036 ( .A(n2325), .B(n3137), .Y(n3550) );
  inv1a1 U4037 ( .A(N661), .Y(n2325) );
  and2a3 U4038 ( .A(N563), .B(n3096), .Y(n3554) );
  and2a3 U4039 ( .A(n3097), .B(reg2[7]), .Y(n3553) );
  and2a3 U4040 ( .A(n3095), .B(reg1[7]), .Y(n3552) );
  and2a3 U4041 ( .A(reg0[7]), .B(n3098), .Y(n3551) );
  inv1a1 U4042 ( .A(n212), .Y(n2402) );
  and2a3 U4043 ( .A(n2996), .B(N947), .Y(n3536) );
  oa1f1 U4044 ( .A(N547), .B(n3143), .C(n3555), .Y(n2323) );
  and2a3 U4045 ( .A(n2624), .B(datai[8]), .Y(n3555) );
  or4a3 U4046 ( .A(n3556), .B(n3557), .C(n3558), .D(n3559), .Y(N5668) );
  or4a3 U4047 ( .A(n3560), .B(n3561), .C(n3562), .D(n3563), .Y(n3559) );
  or3a1 U4048 ( .A(n3564), .B(n3565), .C(n3566), .Y(n3563) );
  and2a3 U4049 ( .A(N1035), .B(n2532), .Y(n3566) );
  and2a3 U4050 ( .A(N2124), .B(n2998), .Y(n3565) );
  and2a3 U4051 ( .A(N3348), .B(n2593), .Y(n3564) );
  and2a3 U4052 ( .A(N2532), .B(n2580), .Y(n3562) );
  and2a3 U4053 ( .A(N3756), .B(n2997), .Y(n3561) );
  and2a3 U4054 ( .A(N2940), .B(n2581), .Y(n3560) );
  or3a1 U4055 ( .A(n3567), .B(n3568), .C(n3569), .Y(n3558) );
  and2a3 U4056 ( .A(N4164), .B(n2582), .Y(n3569) );
  and2a3 U4057 ( .A(N4980), .B(n3000), .Y(n3568) );
  and2a3 U4058 ( .A(N4572), .B(n3001), .Y(n3567) );
  ao1f1 U4059 ( .A(n3159), .B(n2404), .C(n3570), .Y(n3557) );
  or2a1 U4060 ( .A(n2328), .B(n3137), .Y(n3570) );
  inv1a1 U4061 ( .A(N660), .Y(n2328) );
  and2a3 U4062 ( .A(N562), .B(n3096), .Y(n3574) );
  and2a3 U4063 ( .A(n3097), .B(reg2[6]), .Y(n3573) );
  and2a3 U4064 ( .A(n3095), .B(reg1[6]), .Y(n3572) );
  and2a3 U4065 ( .A(reg0[6]), .B(n3098), .Y(n3571) );
  inv1a1 U4066 ( .A(n213), .Y(n2404) );
  and2a3 U4067 ( .A(n2996), .B(N946), .Y(n3556) );
  oa1f1 U4068 ( .A(N548), .B(n3143), .C(n3575), .Y(n2326) );
  and2a3 U4069 ( .A(n2624), .B(datai[7]), .Y(n3575) );
  or4a3 U4070 ( .A(n3576), .B(n3577), .C(n3578), .D(n3579), .Y(N5666) );
  or4a3 U4071 ( .A(n3580), .B(n3581), .C(n3582), .D(n3583), .Y(n3579) );
  or3a1 U4072 ( .A(n3584), .B(n3585), .C(n3586), .Y(n3583) );
  and2a3 U4073 ( .A(N1034), .B(n2532), .Y(n3586) );
  and2a3 U4074 ( .A(N2123), .B(n2998), .Y(n3585) );
  and2a3 U4075 ( .A(N3347), .B(n2593), .Y(n3584) );
  and2a3 U4076 ( .A(N2531), .B(n2580), .Y(n3582) );
  and2a3 U4077 ( .A(N3755), .B(n2997), .Y(n3581) );
  and2a3 U4078 ( .A(N2939), .B(n2581), .Y(n3580) );
  or3a1 U4079 ( .A(n3587), .B(n3588), .C(n3589), .Y(n3578) );
  and2a3 U4080 ( .A(N4163), .B(n2582), .Y(n3589) );
  and2a3 U4081 ( .A(N4979), .B(n3000), .Y(n3588) );
  and2a3 U4082 ( .A(N4571), .B(n3001), .Y(n3587) );
  ao1f1 U4083 ( .A(n3159), .B(n2406), .C(n3590), .Y(n3577) );
  or2a1 U4084 ( .A(n2331), .B(n3137), .Y(n3590) );
  inv1a1 U4085 ( .A(N659), .Y(n2331) );
  and2a3 U4086 ( .A(N561), .B(n3096), .Y(n3594) );
  and2a3 U4087 ( .A(n3097), .B(reg2[5]), .Y(n3593) );
  and2a3 U4088 ( .A(n3095), .B(reg1[5]), .Y(n3592) );
  and2a3 U4089 ( .A(reg0[5]), .B(n3098), .Y(n3591) );
  inv1a1 U4090 ( .A(n214), .Y(n2406) );
  and2a3 U4091 ( .A(n2996), .B(N945), .Y(n3576) );
  oa1f1 U4092 ( .A(N549), .B(n3143), .C(n3595), .Y(n2329) );
  and2a3 U4093 ( .A(n2624), .B(datai[6]), .Y(n3595) );
  or4a3 U4094 ( .A(n3596), .B(n3597), .C(n3598), .D(n3599), .Y(N5664) );
  or4a3 U4095 ( .A(n3600), .B(n3601), .C(n3602), .D(n3603), .Y(n3599) );
  or3a1 U4096 ( .A(n3604), .B(n3605), .C(n3606), .Y(n3603) );
  and2a3 U4097 ( .A(N1033), .B(n2532), .Y(n3606) );
  and2a3 U4098 ( .A(N2122), .B(n2998), .Y(n3605) );
  and2a3 U4099 ( .A(N3346), .B(n2593), .Y(n3604) );
  and2a3 U4100 ( .A(N2530), .B(n2580), .Y(n3602) );
  and2a3 U4101 ( .A(N3754), .B(n2997), .Y(n3601) );
  and2a3 U4102 ( .A(N2938), .B(n2581), .Y(n3600) );
  or3a1 U4103 ( .A(n3607), .B(n3608), .C(n3609), .Y(n3598) );
  and2a3 U4104 ( .A(N4162), .B(n2582), .Y(n3609) );
  and2a3 U4105 ( .A(N4978), .B(n3000), .Y(n3608) );
  and2a3 U4106 ( .A(N4570), .B(n3001), .Y(n3607) );
  ao1f1 U4107 ( .A(n3159), .B(n2408), .C(n3610), .Y(n3597) );
  or2a1 U4108 ( .A(n2334), .B(n3137), .Y(n3610) );
  inv1a1 U4109 ( .A(N658), .Y(n2334) );
  and2a3 U4110 ( .A(N560), .B(n3096), .Y(n3614) );
  and2a3 U4111 ( .A(n3097), .B(reg2[4]), .Y(n3613) );
  and2a3 U4112 ( .A(n3095), .B(reg1[4]), .Y(n3612) );
  and2a3 U4113 ( .A(reg0[4]), .B(n3098), .Y(n3611) );
  inv1a1 U4114 ( .A(n215), .Y(n2408) );
  and2a3 U4115 ( .A(n2996), .B(N944), .Y(n3596) );
  oa1f1 U4116 ( .A(N550), .B(n3143), .C(n3615), .Y(n2332) );
  and2a3 U4117 ( .A(n2624), .B(datai[5]), .Y(n3615) );
  or4a3 U4118 ( .A(n3616), .B(n3617), .C(n3618), .D(n3619), .Y(N5662) );
  or4a3 U4119 ( .A(n3620), .B(n3621), .C(n3622), .D(n3623), .Y(n3619) );
  or3a1 U4120 ( .A(n3624), .B(n3625), .C(n3626), .Y(n3623) );
  and2a3 U4121 ( .A(N1032), .B(n2532), .Y(n3626) );
  and2a3 U4122 ( .A(N2121), .B(n2998), .Y(n3625) );
  and2a3 U4123 ( .A(N3345), .B(n2593), .Y(n3624) );
  and2a3 U4124 ( .A(N2529), .B(n2580), .Y(n3622) );
  and2a3 U4125 ( .A(N3753), .B(n2997), .Y(n3621) );
  and2a3 U4126 ( .A(N2937), .B(n2581), .Y(n3620) );
  or3a1 U4127 ( .A(n3627), .B(n3628), .C(n3629), .Y(n3618) );
  and2a3 U4128 ( .A(N4161), .B(n2582), .Y(n3629) );
  and2a3 U4129 ( .A(N4977), .B(n3000), .Y(n3628) );
  and2a3 U4130 ( .A(N4569), .B(n3001), .Y(n3627) );
  ao1f1 U4131 ( .A(n3159), .B(n2410), .C(n3630), .Y(n3617) );
  or2a1 U4132 ( .A(n2337), .B(n3137), .Y(n3630) );
  inv1a1 U4133 ( .A(N657), .Y(n2337) );
  and2a3 U4134 ( .A(N559), .B(n3096), .Y(n3634) );
  and2a3 U4135 ( .A(reg2[3]), .B(n3097), .Y(n3633) );
  and2a3 U4136 ( .A(reg1[3]), .B(n3095), .Y(n3632) );
  and2a3 U4137 ( .A(reg0[3]), .B(n3098), .Y(n3631) );
  inv1a1 U4138 ( .A(n216), .Y(n2410) );
  and2a3 U4139 ( .A(n2996), .B(N943), .Y(n3616) );
  oa1f1 U4140 ( .A(N551), .B(n3143), .C(n3635), .Y(n2335) );
  and2a3 U4141 ( .A(n2624), .B(datai[4]), .Y(n3635) );
  or4a3 U4142 ( .A(n3636), .B(n3637), .C(n3638), .D(n3639), .Y(N5660) );
  or4a3 U4143 ( .A(n3640), .B(n3641), .C(n3642), .D(n3643), .Y(n3639) );
  or3a1 U4144 ( .A(n3644), .B(n3645), .C(n3646), .Y(n3643) );
  and2a3 U4145 ( .A(N1031), .B(n2532), .Y(n3646) );
  and2a3 U4146 ( .A(N2120), .B(n2998), .Y(n3645) );
  and2a3 U4147 ( .A(N3344), .B(n2593), .Y(n3644) );
  and2a3 U4148 ( .A(N2528), .B(n2580), .Y(n3642) );
  and2a3 U4149 ( .A(N3752), .B(n2997), .Y(n3641) );
  and2a3 U4150 ( .A(N2936), .B(n2581), .Y(n3640) );
  or3a1 U4151 ( .A(n3647), .B(n3648), .C(n3649), .Y(n3638) );
  and2a3 U4152 ( .A(N4160), .B(n2582), .Y(n3649) );
  and2a3 U4153 ( .A(N4976), .B(n3000), .Y(n3648) );
  and2a3 U4154 ( .A(N4568), .B(n3001), .Y(n3647) );
  ao1f1 U4155 ( .A(n3159), .B(n2414), .C(n3650), .Y(n3637) );
  or2a1 U4156 ( .A(n2341), .B(n3137), .Y(n3650) );
  inv1a1 U4157 ( .A(N656), .Y(n2341) );
  and2a3 U4158 ( .A(N558), .B(n3096), .Y(n3654) );
  and2a3 U4159 ( .A(reg2[2]), .B(n3097), .Y(n3653) );
  and2a3 U4160 ( .A(reg1[2]), .B(n3095), .Y(n3652) );
  and2a3 U4161 ( .A(reg0[2]), .B(n3098), .Y(n3651) );
  inv1a1 U4162 ( .A(n217), .Y(n2414) );
  and2a3 U4163 ( .A(n2996), .B(N942), .Y(n3636) );
  oa1f1 U4164 ( .A(N552), .B(n3143), .C(n3655), .Y(n2339) );
  and2a3 U4165 ( .A(n2624), .B(datai[3]), .Y(n3655) );
  or4a3 U4166 ( .A(n3656), .B(n3657), .C(n3658), .D(n3659), .Y(N5658) );
  or4a3 U4167 ( .A(n3660), .B(n3661), .C(n3662), .D(n3663), .Y(n3659) );
  or3a1 U4168 ( .A(n3664), .B(n3665), .C(n3666), .Y(n3663) );
  and2a3 U4169 ( .A(N1030), .B(n2532), .Y(n3666) );
  and2a3 U4170 ( .A(N2119), .B(n2998), .Y(n3665) );
  and2a3 U4171 ( .A(N3343), .B(n2593), .Y(n3664) );
  and2a3 U4172 ( .A(N2527), .B(n2580), .Y(n3662) );
  and2a3 U4173 ( .A(N3751), .B(n2997), .Y(n3661) );
  and2a3 U4174 ( .A(N2935), .B(n2581), .Y(n3660) );
  or3a1 U4175 ( .A(n3667), .B(n3668), .C(n3669), .Y(n3658) );
  and2a3 U4176 ( .A(N4159), .B(n2582), .Y(n3669) );
  and2a3 U4177 ( .A(N4975), .B(n3000), .Y(n3668) );
  and2a3 U4178 ( .A(N4567), .B(n3001), .Y(n3667) );
  ao1f1 U4179 ( .A(n3159), .B(n2436), .C(n3670), .Y(n3657) );
  or2a1 U4180 ( .A(n2364), .B(n3137), .Y(n3670) );
  inv1a1 U4181 ( .A(N655), .Y(n2364) );
  and2a3 U4182 ( .A(N557), .B(n3096), .Y(n3674) );
  and2a3 U4183 ( .A(reg2[1]), .B(n3097), .Y(n3673) );
  and2a3 U4184 ( .A(reg1[1]), .B(n3095), .Y(n3672) );
  and2a3 U4185 ( .A(reg0[1]), .B(n3098), .Y(n3671) );
  inv1a1 U4186 ( .A(n218), .Y(n2436) );
  and2a3 U4187 ( .A(n2996), .B(N941), .Y(n3656) );
  oa1f1 U4188 ( .A(N553), .B(n3143), .C(n3675), .Y(n2362) );
  and2a3 U4189 ( .A(n2624), .B(datai[2]), .Y(n3675) );
  or4a3 U4190 ( .A(n3676), .B(n3677), .C(n3678), .D(n3679), .Y(N5656) );
  or4a3 U4191 ( .A(n3680), .B(n3681), .C(n3682), .D(n3683), .Y(n3679) );
  or3a1 U4192 ( .A(n3684), .B(n3685), .C(n3686), .Y(n3683) );
  and2a3 U4193 ( .A(N1029), .B(n2532), .Y(n3686) );
  and2a3 U4194 ( .A(N2118), .B(n2998), .Y(n3685) );
  and2a3 U4195 ( .A(N3342), .B(n2593), .Y(n3684) );
  and2a3 U4196 ( .A(N2526), .B(n2580), .Y(n3682) );
  and2a3 U4197 ( .A(N3750), .B(n2997), .Y(n3681) );
  and2a3 U4198 ( .A(N2934), .B(n2581), .Y(n3680) );
  or3a1 U4199 ( .A(n3687), .B(n3688), .C(n3689), .Y(n3678) );
  and2a3 U4200 ( .A(N4158), .B(n2582), .Y(n3689) );
  and2a3 U4201 ( .A(N4974), .B(n3000), .Y(n3688) );
  and2a3 U4202 ( .A(N4566), .B(n3001), .Y(n3687) );
  ao1f1 U4203 ( .A(n3159), .B(n2458), .C(n3690), .Y(n3677) );
  or2a1 U4204 ( .A(n2397), .B(n3137), .Y(n3690) );
  inv1a1 U4205 ( .A(n2995), .Y(n2464) );
  inv1a1 U4206 ( .A(N654), .Y(n2397) );
  and2a3 U4207 ( .A(N556), .B(n3096), .Y(n3695) );
  and2a3 U4208 ( .A(reg2[0]), .B(n3097), .Y(n3694) );
  and2a3 U4209 ( .A(reg1[0]), .B(n3095), .Y(n3693) );
  and2a3 U4210 ( .A(reg0[0]), .B(n3098), .Y(n3692) );
  inv1a1 U4211 ( .A(n3696), .Y(n3699) );
  mx2a1 U4212 ( .D0(IR[30]), .D1(n3700), .S(N325), .Y(n3696) );
  xor2a1 U4213 ( .A(N323), .B(n3701), .Y(n3700) );
  and2a3 U4214 ( .A(n3702), .B(n3703), .Y(n3701) );
  inv1a1 U4215 ( .A(n3697), .Y(n3698) );
  xor2a1 U4216 ( .A(n3702), .B(n3703), .Y(n3697) );
  ao1a1 U4217 ( .A(n3704), .B(n3025), .C(n3705), .Y(n3703) );
  or2a1 U4218 ( .A(n3706), .B(n3707), .Y(n3704) );
  mx2a1 U4219 ( .D0(IR[29]), .D1(N322), .S(N325), .Y(n3702) );
  inv1a1 U4220 ( .A(n219), .Y(n2458) );
  and2a3 U4221 ( .A(n2996), .B(N940), .Y(n3676) );
  oa1f1 U4222 ( .A(N554), .B(n3143), .C(n3708), .Y(n2395) );
  and2a3 U4223 ( .A(n2624), .B(datai[1]), .Y(n3708) );
  or4a3 U4224 ( .A(n3709), .B(n3710), .C(n3711), .D(n3712), .Y(N5654) );
  or4a3 U4225 ( .A(n3713), .B(n3714), .C(n3715), .D(n3716), .Y(n3712) );
  or3a1 U4226 ( .A(n3717), .B(n3718), .C(n3719), .Y(n3716) );
  and2a3 U4227 ( .A(N4973), .B(n3000), .Y(n3719) );
  and2a3 U4228 ( .A(N4565), .B(n3001), .Y(n3718) );
  and2a3 U4229 ( .A(n220), .B(n2317), .Y(n3717) );
  and2a3 U4230 ( .A(n3005), .B(n2995), .Y(n2317) );
  and2a3 U4231 ( .A(n3004), .B(n3036), .Y(n2995) );
  or2a1 U4232 ( .A(n3143), .B(n2779), .Y(n3005) );
  and2a3 U4233 ( .A(N3341), .B(n2593), .Y(n3715) );
  and2a3 U4234 ( .A(n2996), .B(N939), .Y(n3714) );
  and2a3 U4235 ( .A(n2624), .B(datai[0]), .Y(n3721) );
  or2a1 U4236 ( .A(n2315), .B(n2316), .Y(n2772) );
  and2a3 U4237 ( .A(n3722), .B(n2755), .Y(n2316) );
  and2a3 U4238 ( .A(n2755), .B(n2756), .Y(n2315) );
  and2a3 U4239 ( .A(n3691), .B(n3722), .Y(n2779) );
  and2a3 U4240 ( .A(n3691), .B(n2756), .Y(n3143) );
  inv1a1 U4241 ( .A(n3722), .Y(n2756) );
  xor2a1 U4242 ( .A(n3705), .B(n3707), .Y(n3722) );
  inv1a1 U4243 ( .A(n2755), .Y(n3691) );
  and2a3 U4244 ( .A(n3707), .B(n3705), .Y(n3723) );
  ao1a1 U4245 ( .A(n3724), .B(n3025), .C(n3021), .Y(n3705) );
  inv1a1 U4246 ( .A(n3725), .Y(n3021) );
  ao1f1 U4247 ( .A(n3026), .B(n3726), .C(n3025), .Y(n3725) );
  or2a1 U4248 ( .A(n3727), .B(n3023), .Y(n3726) );
  mx2a1 U4249 ( .D0(IR[23]), .D1(N316), .S(N325), .Y(n3023) );
  or4a3 U4250 ( .A(n3728), .B(n3729), .C(N536), .D(n3730), .Y(n3026) );
  or3a1 U4251 ( .A(n3020), .B(n3019), .C(n3016), .Y(n3724) );
  mx2a1 U4252 ( .D0(IR[26]), .D1(N319), .S(N325), .Y(n3016) );
  mx2a1 U4253 ( .D0(N318), .D1(IR[25]), .S(n3731), .Y(n3019) );
  mx2a1 U4254 ( .D0(IR[24]), .D1(N317), .S(N325), .Y(n3020) );
  mx2a1 U4255 ( .D0(IR[27]), .D1(N320), .S(N325), .Y(n3707) );
  mx2a1 U4256 ( .D0(IR[28]), .D1(N321), .S(N325), .Y(n3706) );
  and2a3 U4257 ( .A(N4157), .B(n2582), .Y(n3713) );
  and2a3 U4258 ( .A(n3720), .B(n3050), .Y(n3056) );
  or3a1 U4259 ( .A(n3732), .B(n3733), .C(n3734), .Y(n3711) );
  and2a3 U4260 ( .A(N2933), .B(n2581), .Y(n3734) );
  and2a3 U4261 ( .A(N1028), .B(n2532), .Y(n3733) );
  and2a3 U4262 ( .A(N2117), .B(n2998), .Y(n3732) );
  and2a3 U4263 ( .A(N2525), .B(n2580), .Y(n3710) );
  and2a3 U4264 ( .A(N3749), .B(n2997), .Y(n3709) );
  and2a3 U4265 ( .A(n3737), .B(n3728), .Y(n3736) );
  mx2a1 U4266 ( .D0(IR[22]), .D1(N315), .S(N325), .Y(n3729) );
  and2a3 U4267 ( .A(n3730), .B(n3735), .Y(n3737) );
  and2a3 U4268 ( .A(N536), .B(n3027), .Y(n3735) );
  and2a3 U4269 ( .A(n3727), .B(n3025), .Y(n3027) );
  and2a3 U4270 ( .A(N324), .B(N325), .Y(n3025) );
  or4a3 U4271 ( .A(n3738), .B(n3739), .C(n3740), .D(n3741), .Y(n3727) );
  or4a3 U4272 ( .A(n3742), .B(n3743), .C(n3744), .D(n3745), .Y(n3741) );
  or2a1 U4273 ( .A(N552), .B(N551), .Y(n3745) );
  or3a1 U4274 ( .A(N553), .B(N555), .C(N554), .Y(n3744) );
  or2a1 U4275 ( .A(N547), .B(N546), .Y(n3743) );
  or3a1 U4276 ( .A(N548), .B(N550), .C(N549), .Y(n3742) );
  or4a3 U4277 ( .A(N538), .B(N537), .C(N540), .D(N539), .Y(n3740) );
  or2a1 U4278 ( .A(N542), .B(N541), .Y(n3739) );
  or3a1 U4279 ( .A(N543), .B(N545), .C(N544), .Y(n3738) );
  mx2a1 U4280 ( .D0(N313), .D1(IR[20]), .S(n3731), .Y(n3730) );
  mx2a1 U4281 ( .D0(N314), .D1(IR[21]), .S(n3731), .Y(n3728) );
endmodule

